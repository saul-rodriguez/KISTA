VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  LAYER LEF58_TYPE STRING ;
  LAYER LEF58_ENCLOSURE STRING ;
  LAYER LEF58_SPACING STRING ;
  LAYER LEF58_WIDTH STRING ;
  LIBRARY LEF58_MAXVIASTACK STRING "
                        MAXVIASTACK 1 WITHIN Via1 0.99 Via2 0.99 ;" ;
END PROPERTYDEFINITIONS

UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MANUFACTURINGGRID 0.005 ;
LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

LAYER PWdummy
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE PWELL ;" ;
  PROPERTY LEF58_SPACING "SPACING 0.3 ;" ;
  PROPERTY LEF58_WIDTH "WIDTH 0.3 ;" ;
END PWdummy

LAYER Nwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
  PROPERTY LEF58_SPACING "SPACING 0.6 ;
  SPACING 0.24 ;
  SPACING 0.24 ;" ;
  PROPERTY LEF58_WIDTH "WIDTH 0.3 ;" ;
END Nwell

LAYER Oxide
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE DIFFUSION ;" ;
  PROPERTY LEF58_WIDTH "WIDTH 0.05 ;" ;
END Oxide

LAYER Nimp
  TYPE IMPLANT ;
  WIDTH 0.12 ;
  SPACING 0.12 ;
  AREA 0.018 ;
END Nimp

LAYER Pimp
  TYPE IMPLANT ;
  WIDTH 0.12 ;
  SPACING 0.12 ;
  AREA 0.018 ;
END Pimp

LAYER Poly
  TYPE MASTERSLICE ;
END Poly

LAYER Cont
  TYPE CUT ;
  SPACING 0.06 ;
  SPACING 0.08 ADJACENTCUTS 3 WITHIN 0.1 ;
  WIDTH 1 ;
  ENCLOSURE BELOW 0.02 0.03 ;
  ENCLOSURE ABOVE 0 0.03 ;
  DCCURRENTDENSITY AVERAGE 0.1 ;
END Cont

LAYER Metal1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 4 4 ;
  WIDTH 2 ;
  OFFSET 2 2 ;
  SPACING 2 ;
  MINIMUMCUT 2 WIDTH 1.5 FROMABOVE LENGTH 1.5 WITHIN 3 ;
  RESISTANCE RPERSQ 0.0736 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.15 ;
  EDGECAPACITANCE 0.0002 ;
  DCCURRENTDENSITY AVERAGE 2 ;
END Metal1

LAYER Via1
  TYPE CUT ;
  SPACING 1 ;
  WIDTH 1 ;
  ENCLOSURE BELOW 0.005 0.03 ;
  ENCLOSURE ABOVE 0.005 0.03 ;
  RESISTANCE 0.1 ;
  DCCURRENTDENSITY AVERAGE 0.1 ;
END Via1

LAYER Metal2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 4 4 ;
  WIDTH 2 ;
  OFFSET 2 2 ;
  SPACING 2 ;
  MINIMUMCUT 2 WIDTH 1.5 FROMBELOW LENGTH 1.5 WITHIN 3 ;
  MINIMUMCUT 2 WIDTH 1.5 FROMABOVE LENGTH 1.5 WITHIN 3 ;
  RESISTANCE RPERSQ 0.0604 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.18 ;
  EDGECAPACITANCE 0.0002 ;
  DCCURRENTDENSITY AVERAGE 2 ;
END Metal2

LAYER Via2
  TYPE CUT ;
  SPACING 1 ;
  WIDTH 1 ;
  ENCLOSURE BELOW 0.005 0.03 ;
  ENCLOSURE ABOVE 0.005 0.03 ;
  RESISTANCE 0.1 ;
  DCCURRENTDENSITY AVERAGE 0.1 ;
END Via2

LAYER Metal3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 4 4 ;
  WIDTH 2 ;
  OFFSET 2 2 ;
  SPACING 2 ;
  MINIMUMCUT 2 WIDTH 1.5 FROMBELOW LENGTH 1.5 WITHIN 3 ;
  RESISTANCE RPERSQ 0.0604 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.18 ;
  EDGECAPACITANCE 0.0002 ;
  DCCURRENTDENSITY AVERAGE 2 ;
END Metal3

VIARULE M3_M2 GENERATE
  LAYER Metal2 ;
    ENCLOSURE 0.5 0.5 ;
  LAYER Metal3 ;
    ENCLOSURE 0.5 0.5 ;
  LAYER Via2 ;
    RECT -0.5 -0.5 0.5 0.5 ;
    SPACING 2 BY 2 ;
    RESISTANCE 1.000000 ;
END M3_M2

VIARULE M2_M1 GENERATE
  LAYER Metal1 ;
    ENCLOSURE 0.5 0.5 ;
  LAYER Metal2 ;
    ENCLOSURE 0.5 0.5 ;
  LAYER Via1 ;
    RECT -0.5 -0.5 0.5 0.5 ;
    SPACING 2 BY 2 ;
    RESISTANCE 1.000000 ;
END M2_M1

VIARULE M1_PO GENERATE
  LAYER Poly ;
    ENCLOSURE 0.5 0.5 ;
  LAYER Metal1 ;
    ENCLOSURE 0.5 0.5 ;
  LAYER Cont ;
    RECT -0.5 -0.5 0.5 0.5 ;
    SPACING 2 BY 2 ;
    RESISTANCE 1.000000 ;
END M1_PO

VIARULE M1_DIFF GENERATE
  LAYER Oxide ;
    ENCLOSURE 0.5 0.5 ;
  LAYER Metal1 ;
    ENCLOSURE 0.5 0.5 ;
  LAYER Cont ;
    RECT -0.5 -0.5 0.5 0.5 ;
    SPACING 2 BY 2 ;
    RESISTANCE 5.000000 ;
END M1_DIFF

VIARULE M1_PSUB GENERATE
  LAYER Oxide ;
    ENCLOSURE 0.5 0.5 ;
  LAYER Metal1 ;
    ENCLOSURE 0.5 0.5 ;
  LAYER Cont ;
    RECT -0.5 -0.5 0.5 0.5 ;
    SPACING 2 BY 2 ;
    RESISTANCE 5.000000 ;
END M1_PSUB

VIARULE M1_PIMP GENERATE
  LAYER Oxide ;
    ENCLOSURE 0.5 0.5 ;
  LAYER Metal1 ;
    ENCLOSURE 0.5 0.5 ;
  LAYER Cont ;
    RECT -0.5 -0.5 0.5 0.5 ;
    SPACING 2 BY 2 ;
    RESISTANCE 5.000000 ;
END M1_PIMP

VIARULE M1_NIMP GENERATE
  LAYER Oxide ;
    ENCLOSURE 0.5 0.5 ;
  LAYER Metal1 ;
    ENCLOSURE 0.5 0.5 ;
  LAYER Cont ;
    RECT -0.5 -0.5 0.5 0.5 ;
    SPACING 2 BY 2 ;
    RESISTANCE 5.000000 ;
END M1_NIMP

VIARULE M1_NWELL GENERATE
  LAYER Oxide ;
    ENCLOSURE 0.5 0.5 ;
  LAYER Metal1 ;
    ENCLOSURE 0.5 0.5 ;
  LAYER Cont ;
    RECT -0.5 -0.5 0.5 0.5 ;
    SPACING 2 BY 2 ;
    RESISTANCE 5.000000 ;
END M1_NWELL

VIA M2_M1_HV DEFAULT
  LAYER Metal1 ;
    RECT -1 -1 1 1 ;
  LAYER Metal2 ;
    RECT -1 -1 1 1 ;
  LAYER Via1 ;
    RECT -0.5 -0.5 0.5 0.5 ;
END M2_M1_HV

VIA M2_M1_VV DEFAULT
  LAYER Metal1 ;
    RECT -1 -1 1 1 ;
  LAYER Metal2 ;
    RECT -1 -1 1 1 ;
  LAYER Via1 ;
    RECT -0.5 -0.5 0.5 0.5 ;
END M2_M1_VV

VIA M2_M1_VH DEFAULT
  LAYER Metal1 ;
    RECT -1 -1 1 1 ;
  LAYER Metal2 ;
    RECT -1 -1 1 1 ;
  LAYER Via1 ;
    RECT -0.5 -0.5 0.5 0.5 ;
END M2_M1_VH

VIA M2_M1_HH DEFAULT
  LAYER Metal1 ;
    RECT -1 -1 1 1 ;
  LAYER Metal2 ;
    RECT -1 -1 1 1 ;
  LAYER Via1 ;
    RECT -0.5 -0.5 0.5 0.5 ;
END M2_M1_HH

VIA M3_M2_VH DEFAULT
  LAYER Metal2 ;
    RECT -1 -1 1 1 ;
  LAYER Metal3 ;
    RECT -1 -1 1 1 ;
  LAYER Via2 ;
    RECT -0.5 -0.5 0.5 0.5 ;
END M3_M2_VH

VIA M3_M2_HH DEFAULT
  LAYER Metal2 ;
    RECT -1 -1 1 1 ;
  LAYER Metal3 ;
    RECT -1 -1 1 1 ;
  LAYER Via2 ;
    RECT -0.5 -0.5 0.5 0.5 ;
END M3_M2_HH

VIA M3_M2_HV DEFAULT
  LAYER Metal2 ;
    RECT -1 -1 1 1 ;
  LAYER Metal3 ;
    RECT -1 -1 1 1 ;
  LAYER Via2 ;
    RECT -0.5 -0.5 0.5 0.5 ;
END M3_M2_HV

VIA M3_M2_VV DEFAULT
  LAYER Metal2 ;
    RECT -1 -1 1 1 ;
  LAYER Metal3 ;
    RECT -1 -1 1 1 ;
  LAYER Via2 ;
    RECT -0.5 -0.5 0.5 0.5 ;
END M3_M2_VV

NONDEFAULTRULE LEFSpecialRouteSpec
  LAYER Metal1
    WIDTH 2 ;
  END Metal1
  LAYER Metal2
    WIDTH 2 ;
  END Metal2
  LAYER Metal3
    WIDTH 2 ;
  END Metal3
  USEVIARULE M2_M1 ;
  USEVIARULE M3_M2 ;
END LEFSpecialRouteSpec
NONDEFAULTRULE VLMDefaultSetup
  LAYER Metal1
    WIDTH 2 ;
  END Metal1
  LAYER Metal2
    WIDTH 2 ;
  END Metal2
  LAYER Metal3
    WIDTH 2 ;
  END Metal3
  USEVIARULE M1_PO ;
  USEVIARULE M1_NWELL ;
  USEVIARULE M1_PSUB ;
  USEVIARULE M1_NIMP ;
  USEVIARULE M1_PIMP ;
  USEVIARULE M1_DIFF ;
  USEVIARULE M2_M1 ;
  USEVIARULE M3_M2 ;
END VLMDefaultSetup
SITE CoreSite
  CLASS CORE ;
  SIZE 4 BY 40 ;
END CoreSite

SITE IOSite
  CLASS PAD ;
  SIZE 1 BY 240 ;
END IOSite

SITE CornerSite
  CLASS PAD ;
  SIZE 240 BY 240 ;
END CornerSite

SITE CoreSiteDouble
  CLASS CORE ;
  SIZE 4 BY 80 ;
END CoreSiteDouble

END LIBRARY
