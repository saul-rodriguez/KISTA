//Verilog HDL for "KISTA_SOI_STDLIB2", "TIELO" "functional"


`timescale 1ns/10ps
`celldefine
module TIELO (Y);
	output Y;
	//input A;

	// Function
	buf (Y, 1'b0);

	// Timing
	specify
	endspecify
endmodule
`endcelldefine
