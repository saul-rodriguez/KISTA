*
*
*
*                       LINUX           Tue Dec 21 07:14:31 2021
*
*
*
*  PROGRAM  advgen
*
*  Name           : advgen - Quantus - (64-bit)
*  Version        : 20.1.2-p025
*  Build Date     : Thu Sep 3 13:54:09 PDT 2020
*
*  HSPICE LIBRARY
*
*
*

*
.GLOBAL VSS! VDD!
.SUBCKT OAI21X1 B0 Y A0 A1
*
*
*  caps2d version: 10
*
*
*       TRANSISTOR CARDS
*
*
MX5_M0_unmatched	Y#3	B0#6	net13#4	net13#4	nch
+ L=1e-06	W=4e-06
+ AD=1e-11	AS=0	PD=1.3e-05	PS=0
+ fw=4e-06 sa=2e-06 sb=2e-06
MX4_M0_unmatched	net13#2	A1#4	VSS!#3	VSS!#3	nch	L=1e-06
+ W=4e-06
+ AD=1e-11	AS=0	PD=1.3e-05	PS=0
+ fw=4e-06 sa=2e-06 sb=2e-06
MX3_M0_unmatched	net13	A0#4	VSS!#1	VSS!#1	nch	L=1e-06
+ W=4e-06
+ AD=1e-11	AS=0	PD=1.3e-05	PS=0
+ fw=4e-06 sa=2e-06 sb=2e-06
MX8_M0_unmatched	Y#4	B0#4	VDD!#1	VDD!#1	pch	L=1e-06
+ W=8e-06
+ AD=2e-11	AS=0	PD=2.1e-05	PS=0
+ fw=8e-06 sa=2e-06 sb=2e-06
MX7_M0_unmatched	Y#2	A1#2	net15	net15	pch	L=1e-06
+ W=8e-06
+ AD=2e-11	AS=0	PD=2.1e-05	PS=0
+ fw=8e-06 sa=2e-06 sb=2e-06
MX6_M0_unmatched	net15#2	A0#2	VDD!#2	VDD!#2	pch	L=1e-06
+ W=8e-06
+ AD=2e-11	AS=0	PD=2.1e-05	PS=0
+ fw=8e-06 sa=2e-06 sb=2e-06
*
*
*       RESISTOR AND CAP/DIODE CARDS
*
Rd7	B0#4	B0#5	 1636.0317
Rd9	B0#5	B0	   85.4740
Rd8	Y	Y#4	    2.2262
Rd1	Y	Y#2	    2.3261
Rd3	A0#3	A0#4	 2236.0317
Rd2	A1#2	A1#3	 1036.0317
Rd4	A1#3	A1	   85.4640
Rd6	net13#4	net13	    8.7045
Rd5	VSS!	VSS!#3	    3.0612
Rc4	B0#5	B0#6	 1036.0317
Rc14	VDD!#1	VDD!	    1.8054	$metal1_conn
Rc15	VDD!	VDD!#2	    1.5019	$metal1_conn
Rc2	net15	net15#2	    2.7059	$metal1_conn
Rc5	Y	Y#3	    2.6175
Rc6	Y#4	Y#2	    6.6694
Rc12	A0#2	A0#3	  436.0318
Rc10	A0#3	A0	   85.4740
Rc13	A1#3	A1#4	 1636.0317
Rc11	net13#4	net13#2	    7.2395
Rc1	net13#2	net13	    8.4101
Rc3	VSS!#3	VSS!#1	   31.9527
Rc8	VSS!	VSS!#1	    2.9720
Rs1	4	VSS!	50

*
*       CAPACITOR CARDS
*
*
C1	Y	B0	4.0945e-16
C2	B0#4	Y	8.63743e-16
C3	Y#3	B0#6	2.23289e-16
C4	VSS!	B0	1.25563e-17
C5	B0#4	VSS!	6.24104e-18
C6	VSS!#1	B0#6	6.51585e-17
C7	VDD!#1	B0#4	3.44382e-16
C8	4	B0	4.91506e-15
C9	B0#4	4	1.43864e-15
C10	B0#6	4	1.44686e-15
C11	B0#5	4	5.57378e-19
C12	net13#4	B0	6.79721e-18
C13	net13#4	B0#6	1.46232e-16
C14	net13#2	B0	5.50113e-18
C15	B0#4	X8_5	5.0867e-16
C16	VSS!	Y	1.77406e-17
C17	VSS!#1	Y#3	6.81642e-17
C18	Y#4	VDD!#1	2.51355e-16
C19	Y#2	VDD!	6.36186e-17
C20	A1	Y	9.80229e-18
C21	Y#2	A1#2	2.57023e-16
C22	A1#3	Y	6.09111e-19
C23	4	Y	4.68705e-15
C24	Y#3	4	5.35387e-16
C25	net13#4	Y#3	7.91422e-17
C26	net13#2	Y	1.71811e-17
C27	Y#2	net15	1.4059e-16
C28	X8_5	Y	3.32712e-16
C29	X7_5	Y	7.9727e-17
C30	Y#2	X7_5	8.80485e-17
C31	VSS!	A0	1.74085e-17
C32	A0#2	VSS!	2.33242e-18
C33	VSS!#1	A0#4	2.26587e-16
C34	A0#3	VSS!	6.18207e-19
C35	VDD!#2	A0	5.77159e-17
C36	VDD!#2	A0#2	3.4549e-16
C37	A0#3	VDD!#2	7.41669e-19
C38	4	A0	4.76614e-15
C39	A0#2	4	2.60449e-16
C40	A0#4	4	2.62846e-15
C41	A0#3	4	2.73703e-16
C42	A0#4	net13	7.79727e-16
C43	net15#2	A0#2	2.48735e-16
C44	A0#2	X6_5	5.03676e-16
C45	VDD!#2	VSS!	6.38307e-18
C46	A1	VSS!	1.89117e-17
C47	A1#2	VSS!	7.24756e-18
C48	VSS!#3	A1#4	2.11778e-16
C49	A1#3	VSS!	1.17516e-18
C50	4	VSS!	1.26675e-15
C51	VSS!#3	4	2.25171e-16
C52	VSS!#1	4	5.44375e-15
C53	VSS!#3	net13#2	2.06715e-16
C54	VSS!#1	net13	2.78956e-16
C55	net15#2	VSS!	5.05691e-18
C56	A1#2	VDD!	6.39776e-17
C57	4	VDD!	2.55705e-15
C58	VDD!#1	4	2.69303e-15
C59	VDD!#2	4	1.27811e-15
C60	net15	VDD!	7.20445e-17
C61	net15#2	VDD!	6.41265e-17
C62	VDD!#2	net15#2	1.39862e-16
C63	VDD!#1	X8_5	6.48336e-16
C64	X7_5	VDD!	2.866e-17
C65	X6_5	VDD!	2.866e-17
C66	VDD!#2	X6_5	6.48336e-16
C67	4	A1	4.95189e-15
C68	A1#2	4	9.7449e-16
C69	A1#4	4	1.95581e-15
C70	A1#3	4	3.07708e-16
C71	net13#2	A1	1.16618e-17
C72	net13#2	A1#4	7.92435e-16
C73	A1#3	net13#2	7.24662e-19
C74	net15	A1	1.10458e-17
C75	A1#2	net15	2.47812e-16
C76	A1#3	net15	6.86382e-19
C77	A1#2	X7_5	5.22291e-16
C78	net13	4	2.23486e-15
C79	net13#4	4	2.9116e-16
C80	net13#2	4	1.74972e-15
C81	net15	4	1.12243e-16
C82	net15#2	4	5.01172e-17
C83	X7_5	net15	1.78573e-16
C84	net15#2	X6_5	1.7863e-16
*
*
.ENDS OAI21X1
*
