//Verilog HDL for "KISTA_SOI_STDLIB", "DECAP4" "functional"


module DECAP4 ( );

endmodule
