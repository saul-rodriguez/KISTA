//Verilog HDL for "KISTA_SOI_STDLIB", "DECAP2" "functional"


module DECAP2 ( );

endmodule
