//Verilog HDL for "KISTA_SOI_STDLIB2", "AND2X1" "functional"


module AND2X1 (A, B, Y);
	input A, B;
	output Y;

	assign Y = A & B;

endmodule
