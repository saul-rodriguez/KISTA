//Verilog HDL for "KISTA_SOI_STDLIB2", "OR2X1" "functional"


module OR2X1 (A, B, Y, YN );
	input A, B;
	output Y, YN;

	assign Y = A | B;
	assign YN = ~(A | B);

endmodule
