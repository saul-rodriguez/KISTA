//Verilog HDL for "KISTA_SOI_STDLIB", "TIEHI" "functional"


`timescale 1ns/10ps
`celldefine
module TIEHI (Y);
	output Y;


	// Function
	buf (Y, 1'b1);

	// Timing
	specify
	endspecify
endmodule
`endcelldefine