*
*
*
*                       LINUX           Tue Dec 21 14:10:17 2021
*
*
*
*  PROGRAM  advgen
*
*  Name           : advgen - Quantus - (64-bit)
*  Version        : 20.1.2-p025
*  Build Date     : Thu Sep 3 13:54:09 PDT 2020
*
*  HSPICE LIBRARY
*
*
*

*
.GLOBAL VDD! VSS! 
.SUBCKT NOR3X1 Y C A B
*
*
*  caps2d version: 10
*
*
*       TRANSISTOR CARDS
*
*
MX5_M0_unmatched	Y#5	C#4	VSS!#1	VSS!#1	nch	L=1e-06
+ W=2e-06
+ AD=5e-12	AS=0	PD=9e-06	PS=0
+ fw=2e-06 sa=2e-06 sb=2e-06
MX4_M0_unmatched	Y#6	B#4	VSS!#4	VSS!#4	nch	L=1e-06
+ W=2e-06
+ AD=5e-12	AS=0	PD=9e-06	PS=0
+ fw=2e-06 sa=2e-06 sb=2e-06
MX3_M0_unmatched	Y#3	A#4	VSS!#3	VSS!#3	nch	L=1e-06
+ W=2e-06
+ AD=5e-12	AS=0	PD=9e-06	PS=0
+ fw=2e-06 sa=2e-06 sb=2e-06
MX8_M0_unmatched	Y#4	C#2	net60	net60	pch	L=1e-06
+ W=1.2e-05
+ AD=3e-11	AS=0	PD=2.9e-05	PS=0
+ fw=1.2e-05 sa=2e-06 sb=2e-06
MX7_M0_unmatched	net60#2	B#2	net61	net61	pch	L=1e-06
+ W=1.2e-05
+ AD=3e-11	AS=0	PD=2.9e-05	PS=0
+ fw=1.2e-05 sa=2e-06 sb=2e-06
MX6_M0_unmatched	net61#2	A#2	VDD!#1	VDD!#1	pch	L=1e-06
+ W=1.2e-05
+ AD=3e-11	AS=0	PD=2.9e-05	PS=0
+ fw=1.2e-05 sa=2e-06 sb=2e-06
*
*
*       RESISTOR AND CAP/DIODE CARDS
*
Rd7	C#2	C#3	  436.0318
Rd9	C#3	C	   85.4715
Rd8	A#3	A#4	  736.0318
Rd1	VSS!	VSS!#3	    5.2019
Rd3	VSS!#1	VSS!#4	  364.9153
Rd2	B#2	B#3	 1036.0317
Rd4	B#3	B	   85.4690
Rd6	Y	Y#5	    6.3778
Rd5	Y#5	Y#2	   26.2936
Rc16	VDD!	VDD!#1	    1.0827	$metal1_conn
Rc2	net61	net61#2	    1.9725	$metal1_conn
Rc4	net60	net60#2	    1.9725	$metal1_conn
Rc9	C#3	C#4	 1936.0317
Rc6	A#2	A#3	 1636.0317
Rc10	A#3	A	   85.4640
Rc11	VSS!	VSS!#1	    5.4301
Rc8	VSS!	VSS!#4	    5.2279
Rc7	B#3	B#4	 1336.0317
Rc5	Y	Y#4	    1.2633
Rc1	Y	Y#2	    0.2222
Rc14	Y#2	Y#6	    5.0795
Rc13	Y#2	Y#3	    5.2760
Rs1	4	VSS!	50
*
*       CAPACITOR CARDS
*
*
C1	C#4	Y	7.79045e-16
C2	Y#4	C	3.64655e-16
C3	Y#4	C#2	3.72194e-16
C4	Y#4	VDD!	6.62687e-17
C5	Y#3	A	9.04369e-17
C6	Y#3	A#4	1.36031e-16
C7	A#3	Y#3	5.61971e-18
C8	VSS!#1	Y#5	1.26646e-16
C9	Y#3	VSS!	2.37408e-16
C10	Y#2	VSS!#4	8.01849e-17
C11	Y#2	B	2.72725e-17
C12	Y#2	B#4	7.27572e-16
C13	Y#2	B#3	1.6964e-18
C14	4	Y	7.48094e-15
C15	Y#4	net60	2.1454e-16
C16	Y#2	net60#2	2.85752e-18
C17	Y#4	X8_5	8.34381e-16
C18	C#2	VDD!	6.39776e-17
C19	VSS!	C	1.5276e-17
C20	C#2	VSS!	3.29873e-18
C21	VSS!#1	C#4	1.79769e-16
C22	4	C	4.44111e-15
C23	C#2	4	2.58954e-16
C24	C#4	4	2.29314e-15
C25	C#3	4	3.68858e-19
C26	net60	C	5.21191e-17
C27	C#2	net60	3.57573e-16
C28	C#2	X8_5	5.26341e-16
C29	VDD!#1	A#2	4.53526e-16
C30	VDD!#1	VSS!	1.553e-17
C31	B#2	VDD!	6.39776e-17
C32	4	VDD!	6.09126e-15
C33	VDD!#1	4	2.94187e-16
C34	net61	VDD!	7.29903e-17
C35	net61#2	VDD!	6.48416e-17
C36	VDD!#1	net61#2	2.07561e-16
C37	net60	VDD!	1.49785e-16
C38	X7_5	VDD!	2.866e-17
C39	X6_5	VDD!	3.4392e-17
C40	VDD!#1	X6_5	8.34381e-16
C41	VSS!	A	1.64815e-17
C42	A#2	VSS!	3.66463e-18
C43	VSS!#3	A	2.39434e-17
C44	VSS!#3	A#4	1.89046e-16
C45	A#3	VSS!	1.04732e-18
C46	4	A	4.36069e-15
C47	A#2	4	1.67969e-15
C48	A#4	4	1.13196e-15
C49	A#3	4	2.49118e-16
C50	net61#2	A#2	3.58496e-16
C51	A#2	X6_5	5.02932e-16
C52	B	VSS!	1.57514e-17
C53	B#2	VSS!	1.18177e-17
C54	VSS!#4	B#4	1.83665e-16
C55	B#3	VSS!	9.79766e-19
C56	4	VSS!	2.78463e-15
C57	VSS!#1	4	2.76743e-15
C58	VSS!#4	4	1.86083e-16
C59	VSS!#3	4	1.67976e-15
C60	net61	VSS!	6.01843e-18
C61	net60#2	VSS!	2.94747e-18
C62	X8_5	VSS!	5.732e-18
C63	4	B	4.68969e-15
C64	B#2	4	9.39673e-16
C65	B#4	4	1.68242e-15
C66	B#3	4	2.91707e-16
C67	net61	B	1.16185e-17
C68	B#2	net61	3.57573e-16
C69	B#3	net61	7.22692e-19
C70	net60#2	B#2	3.58496e-16
C71	B#2	X7_5	5.22396e-16
C72	net61	4	1.62667e-16
C73	net60#2	4	1.00044e-16
C74	net60#2	net61	2.08289e-16
C75	X7_5	net61	1.78672e-16
C76	net61#2	X6_5	1.78672e-16
C77	X8_5	net60	1.78672e-16
C78	net60#2	X7_5	1.78672e-16
*
*
.ENDS NOR3X1
*
