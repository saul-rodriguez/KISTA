//Verilog HDL for "KISTA_SOI_STDLIB2", "NAND2X1" "functional"

// type:  
`timescale 1ns/10ps
`celldefine
module NAND2X3 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire int_fwire_0;

	and (int_fwire_0, A, B);
	not (Y, int_fwire_0);

	// Timing
	specify
		(A => Y) = 0;
		(B => Y) = 0;
	endspecify
endmodule
`endcelldefine