//Verilog HDL for "KISTA_SOI_STDLIB", "DECAP1" "functional"


module DECAP1 ( );

endmodule
