//Verilog HDL for "KISTA_SOI_STDLIB2", "INVX1" "functional"


`timescale 1ns/10ps
`celldefine
module INVX3 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		(A => Y) = 0;
	endspecify
endmodule
`endcelldefine