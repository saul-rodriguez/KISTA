//Verilog HDL for "KISTA_SOI_STDLIB2", "DECAP2" "functional"


module DECAP2 ( );

endmodule
