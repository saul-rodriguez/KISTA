VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO ADDFX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFX1 0 0 ;
  SIZE 124 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 124 3 ;
        RECT 117 -3 119 7 ;
        RECT 97 -3 99 7 ;
        RECT 89 -3 91 7 ;
        RECT 81 -3 83 7 ;
        RECT 73 -3 75 7 ;
        RECT 37 9 47 11 ;
        RECT 45 -3 47 11 ;
        RECT 1 9 15 11 ;
        RECT 1 -3 3 11 ;
    END
  END VSS!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 124 43 ;
        RECT 117 31 119 43 ;
        RECT 87 33 91 43 ;
        RECT 79 33 83 43 ;
        RECT 71 33 75 43 ;
        RECT 45 29 47 43 ;
        RECT 37 29 47 31 ;
        RECT 1 29 9 31 ;
        RECT 1 29 3 43 ;
    END
  END VDD!
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5 17 103 19 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9 13 95 15 ;
    END
  END A
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 121 5 123 35 ;
    END
  END SUM
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 17 21 111 23 ;
    END
  END CIN
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 49 5 71 7 ;
        RECT 49 5 51 11 ;
    END
  END COUT
  OBS
    LAYER Metal1 ;
      RECT 113 5 115 35 ;
      RECT 61 25 63 33 ;
      RECT 57 25 119 27 ;
      RECT 109 29 111 35 ;
      RECT 103 29 111 31 ;
      RECT 65 29 67 33 ;
      RECT 65 29 99 31 ;
      RECT 29 25 33 31 ;
      RECT 21 25 47 27 ;
      RECT 105 5 111 7 ;
      RECT 97 9 107 11 ;
      RECT 95 33 107 35 ;
      RECT 65 9 91 11 ;
      RECT 57 9 63 11 ;
      RECT 49 31 55 35 ;
      RECT 5 33 41 35 ;
      RECT 29 5 39 7 ;
      RECT 21 9 35 11 ;
      RECT 13 29 25 31 ;
      RECT 5 5 23 7 ;
    LAYER Via1 ;
      RECT 121.5 5.5 122.5 6.5 ;
      RECT 121.5 31.5 122.5 32.5 ;
      RECT 121.5 33.5 122.5 34.5 ;
      RECT 117.5 5.5 118.5 6.5 ;
      RECT 117.5 25.5 118.5 26.5 ;
      RECT 117.5 31.5 118.5 32.5 ;
      RECT 117.5 33.5 118.5 34.5 ;
      RECT 113.5 5.5 114.5 6.5 ;
      RECT 113.5 31.5 114.5 32.5 ;
      RECT 113.5 33.5 114.5 34.5 ;
      RECT 109.5 5.5 110.5 6.5 ;
      RECT 109.5 21.5 110.5 22.5 ;
      RECT 109.5 31.5 110.5 32.5 ;
      RECT 109.5 33.5 110.5 34.5 ;
      RECT 105.5 5.5 106.5 6.5 ;
      RECT 105.5 9.5 106.5 10.5 ;
      RECT 105.5 29.5 106.5 30.5 ;
      RECT 105.5 33.5 106.5 34.5 ;
      RECT 103.5 29.5 104.5 30.5 ;
      RECT 103.5 33.5 104.5 34.5 ;
      RECT 101.5 17.5 102.5 18.5 ;
      RECT 97.5 5.5 98.5 6.5 ;
      RECT 97.5 9.5 98.5 10.5 ;
      RECT 97.5 29.5 98.5 30.5 ;
      RECT 97.5 33.5 98.5 34.5 ;
      RECT 95.5 29.5 96.5 30.5 ;
      RECT 95.5 33.5 96.5 34.5 ;
      RECT 93.5 13.5 94.5 14.5 ;
      RECT 89.5 5.5 90.5 6.5 ;
      RECT 89.5 9.5 90.5 10.5 ;
      RECT 89.5 29.5 90.5 30.5 ;
      RECT 89.5 33.5 90.5 34.5 ;
      RECT 87.5 29.5 88.5 30.5 ;
      RECT 87.5 33.5 88.5 34.5 ;
      RECT 85.5 21.5 86.5 22.5 ;
      RECT 81.5 5.5 82.5 6.5 ;
      RECT 81.5 9.5 82.5 10.5 ;
      RECT 81.5 29.5 82.5 30.5 ;
      RECT 81.5 33.5 82.5 34.5 ;
      RECT 79.5 29.5 80.5 30.5 ;
      RECT 79.5 33.5 80.5 34.5 ;
      RECT 77.5 17.5 78.5 18.5 ;
      RECT 73.5 5.5 74.5 6.5 ;
      RECT 73.5 9.5 74.5 10.5 ;
      RECT 73.5 29.5 74.5 30.5 ;
      RECT 73.5 33.5 74.5 34.5 ;
      RECT 71.5 29.5 72.5 30.5 ;
      RECT 71.5 33.5 72.5 34.5 ;
      RECT 69.5 13.5 70.5 14.5 ;
      RECT 65.5 9.5 66.5 10.5 ;
      RECT 65.5 29.5 66.5 30.5 ;
      RECT 65.5 31.5 66.5 32.5 ;
      RECT 61.5 9.5 62.5 10.5 ;
      RECT 61.5 29.5 62.5 30.5 ;
      RECT 61.5 31.5 62.5 32.5 ;
      RECT 57.5 9.5 58.5 10.5 ;
      RECT 57.5 25.5 58.5 26.5 ;
      RECT 53.5 5.5 54.5 6.5 ;
      RECT 53.5 31.5 54.5 32.5 ;
      RECT 53.5 33.5 54.5 34.5 ;
      RECT 49.5 5.5 50.5 6.5 ;
      RECT 49.5 31.5 50.5 32.5 ;
      RECT 49.5 33.5 50.5 34.5 ;
      RECT 45.5 5.5 46.5 6.5 ;
      RECT 45.5 25.5 46.5 26.5 ;
      RECT 45.5 31.5 46.5 32.5 ;
      RECT 45.5 33.5 46.5 34.5 ;
      RECT 43.5 13.5 44.5 14.5 ;
      RECT 39.5 29.5 40.5 30.5 ;
      RECT 39.5 33.5 40.5 34.5 ;
      RECT 37.5 5.5 38.5 6.5 ;
      RECT 37.5 9.5 38.5 10.5 ;
      RECT 37.5 29.5 38.5 30.5 ;
      RECT 37.5 33.5 38.5 34.5 ;
      RECT 33.5 9.5 34.5 10.5 ;
      RECT 33.5 25.5 34.5 26.5 ;
      RECT 31.5 29.5 32.5 30.5 ;
      RECT 31.5 33.5 32.5 34.5 ;
      RECT 29.5 5.5 30.5 6.5 ;
      RECT 29.5 9.5 30.5 10.5 ;
      RECT 29.5 29.5 30.5 30.5 ;
      RECT 29.5 33.5 30.5 34.5 ;
      RECT 25.5 17.5 26.5 18.5 ;
      RECT 25.5 21.5 26.5 22.5 ;
      RECT 23.5 25.5 24.5 26.5 ;
      RECT 23.5 29.5 24.5 30.5 ;
      RECT 21.5 5.5 22.5 6.5 ;
      RECT 21.5 9.5 22.5 10.5 ;
      RECT 21.5 25.5 22.5 26.5 ;
      RECT 21.5 29.5 22.5 30.5 ;
      RECT 17.5 21.5 18.5 22.5 ;
      RECT 15.5 29.5 16.5 30.5 ;
      RECT 15.5 33.5 16.5 34.5 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 9.5 14.5 10.5 ;
      RECT 13.5 29.5 14.5 30.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 13.5 10.5 14.5 ;
      RECT 7.5 29.5 8.5 30.5 ;
      RECT 7.5 33.5 8.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 9.5 6.5 10.5 ;
      RECT 5.5 17.5 6.5 18.5 ;
      RECT 5.5 29.5 6.5 30.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
  END
END ADDFX1

MACRO ADDHX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDHX1 0 0 ;
  SIZE 56 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 56 3 ;
        RECT 49 -3 51 11 ;
        RECT 45 -3 47 11 ;
        RECT 33 -3 35 11 ;
        RECT 17 -3 19 11 ;
        RECT 1 -3 3 11 ;
    END
  END VSS!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 56 43 ;
        RECT 49 27 51 43 ;
        RECT 33 27 35 43 ;
        RECT 29 27 31 43 ;
        RECT 17 27 19 43 ;
        RECT 13 27 15 43 ;
        RECT 1 27 3 43 ;
    END
  END VDD!
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 21 9 23 31 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 53 9 55 31 ;
    END
  END SUM
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5 13 11 15 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 17 3 23 ;
    END
  END A
  OBS
    LAYER Metal1 ;
      RECT 45 17 47 31 ;
      RECT 25 9 27 31 ;
      RECT 25 17 51 19 ;
      RECT 29 13 43 15 ;
      RECT 41 9 43 15 ;
      RECT 37 9 39 15 ;
      RECT 29 9 31 15 ;
      RECT 5 27 11 31 ;
      RECT 9 17 11 31 ;
      RECT 9 17 19 19 ;
      RECT 13 9 15 19 ;
      RECT 37 27 43 31 ;
      RECT 5 9 11 11 ;
    LAYER Via1 ;
      RECT 53.5 9.5 54.5 10.5 ;
      RECT 53.5 27.5 54.5 28.5 ;
      RECT 53.5 29.5 54.5 30.5 ;
      RECT 49.5 9.5 50.5 10.5 ;
      RECT 49.5 17.5 50.5 18.5 ;
      RECT 49.5 27.5 50.5 28.5 ;
      RECT 49.5 29.5 50.5 30.5 ;
      RECT 45.5 9.5 46.5 10.5 ;
      RECT 45.5 27.5 46.5 28.5 ;
      RECT 45.5 29.5 46.5 30.5 ;
      RECT 41.5 9.5 42.5 10.5 ;
      RECT 41.5 27.5 42.5 28.5 ;
      RECT 41.5 29.5 42.5 30.5 ;
      RECT 37.5 9.5 38.5 10.5 ;
      RECT 37.5 27.5 38.5 28.5 ;
      RECT 37.5 29.5 38.5 30.5 ;
      RECT 33.5 9.5 34.5 10.5 ;
      RECT 33.5 27.5 34.5 28.5 ;
      RECT 33.5 29.5 34.5 30.5 ;
      RECT 29.5 9.5 30.5 10.5 ;
      RECT 29.5 27.5 30.5 28.5 ;
      RECT 29.5 29.5 30.5 30.5 ;
      RECT 25.5 9.5 26.5 10.5 ;
      RECT 25.5 27.5 26.5 28.5 ;
      RECT 25.5 29.5 26.5 30.5 ;
      RECT 21.5 9.5 22.5 10.5 ;
      RECT 21.5 27.5 22.5 28.5 ;
      RECT 21.5 29.5 22.5 30.5 ;
      RECT 17.5 9.5 18.5 10.5 ;
      RECT 17.5 17.5 18.5 18.5 ;
      RECT 17.5 27.5 18.5 28.5 ;
      RECT 17.5 29.5 18.5 30.5 ;
      RECT 13.5 9.5 14.5 10.5 ;
      RECT 13.5 27.5 14.5 28.5 ;
      RECT 13.5 29.5 14.5 30.5 ;
      RECT 9.5 9.5 10.5 10.5 ;
      RECT 9.5 13.5 10.5 14.5 ;
      RECT 9.5 27.5 10.5 28.5 ;
      RECT 9.5 29.5 10.5 30.5 ;
      RECT 5.5 9.5 6.5 10.5 ;
      RECT 5.5 27.5 6.5 28.5 ;
      RECT 5.5 29.5 6.5 30.5 ;
      RECT 1.5 9.5 2.5 10.5 ;
      RECT 1.5 17.5 2.5 18.5 ;
      RECT 1.5 27.5 2.5 28.5 ;
      RECT 1.5 29.5 2.5 30.5 ;
  END
END ADDHX1

MACRO AND2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X1 0 0 ;
  SIZE 24 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN YN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5 25 19 27 ;
        RECT 13 5 15 35 ;
        RECT 5 25 7 35 ;
    END
  END YN
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 24 43 ;
        RECT 17 31 19 43 ;
        RECT 9 31 11 43 ;
        RECT 1 31 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 21 3 27 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9 13 11 19 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 21 5 23 35 ;
    END
  END Y
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 24 3 ;
        RECT 17 -3 19 7 ;
        RECT 1 -3 3 7 ;
    END
  END VSS!
  OBS
    LAYER Metal1 ;
      RECT 5 5 11 7 ;
    LAYER Via1 ;
      RECT 21.5 5.5 22.5 6.5 ;
      RECT 21.5 31.5 22.5 32.5 ;
      RECT 21.5 33.5 22.5 34.5 ;
      RECT 17.5 5.5 18.5 6.5 ;
      RECT 17.5 25.5 18.5 26.5 ;
      RECT 17.5 31.5 18.5 32.5 ;
      RECT 17.5 33.5 18.5 34.5 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 13.5 10.5 14.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 21.5 2.5 22.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END AND2X1

MACRO AND3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3X1 0 0 ;
  SIZE 32 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN YN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5 25 27 27 ;
        RECT 21 5 23 35 ;
        RECT 13 25 15 35 ;
        RECT 5 25 7 35 ;
    END
  END YN
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 32 43 ;
        RECT 25 31 27 43 ;
        RECT 17 31 19 43 ;
        RECT 9 31 11 43 ;
        RECT 1 31 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 21 3 27 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9 13 11 19 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 17 9 19 15 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 29 5 31 35 ;
    END
  END Y
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 32 3 ;
        RECT 25 -3 27 7 ;
        RECT 1 -3 3 7 ;
    END
  END VSS!
  OBS
    LAYER Metal1 ;
      RECT 13 5 19 7 ;
      RECT 5 5 11 7 ;
    LAYER Via1 ;
      RECT 29.5 5.5 30.5 6.5 ;
      RECT 29.5 31.5 30.5 32.5 ;
      RECT 29.5 33.5 30.5 34.5 ;
      RECT 25.5 5.5 26.5 6.5 ;
      RECT 25.5 25.5 26.5 26.5 ;
      RECT 25.5 31.5 26.5 32.5 ;
      RECT 25.5 33.5 26.5 34.5 ;
      RECT 21.5 5.5 22.5 6.5 ;
      RECT 21.5 31.5 22.5 32.5 ;
      RECT 21.5 33.5 22.5 34.5 ;
      RECT 17.5 5.5 18.5 6.5 ;
      RECT 17.5 13.5 18.5 14.5 ;
      RECT 17.5 31.5 18.5 32.5 ;
      RECT 17.5 33.5 18.5 34.5 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 13.5 10.5 14.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 21.5 2.5 22.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END AND3X1

MACRO AND4X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4X1 0 0 ;
  SIZE 40 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN YN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5 25 35 27 ;
        RECT 29 5 31 35 ;
        RECT 21 25 23 35 ;
        RECT 13 25 15 35 ;
        RECT 5 25 7 35 ;
    END
  END YN
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 40 43 ;
        RECT 33 31 35 43 ;
        RECT 25 31 27 43 ;
        RECT 17 31 19 43 ;
        RECT 9 31 11 43 ;
        RECT 1 31 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 21 3 27 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9 17 15 19 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 17 13 19 19 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 25 9 27 15 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 37 5 39 35 ;
    END
  END Y
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 40 3 ;
        RECT 33 -3 35 7 ;
        RECT 1 -3 3 7 ;
    END
  END VSS!
  OBS
    LAYER Metal1 ;
      RECT 21 5 27 7 ;
      RECT 13 5 19 7 ;
      RECT 5 5 11 7 ;
    LAYER Via1 ;
      RECT 37.5 5.5 38.5 6.5 ;
      RECT 37.5 31.5 38.5 32.5 ;
      RECT 37.5 33.5 38.5 34.5 ;
      RECT 33.5 5.5 34.5 6.5 ;
      RECT 33.5 25.5 34.5 26.5 ;
      RECT 33.5 31.5 34.5 32.5 ;
      RECT 33.5 33.5 34.5 34.5 ;
      RECT 29.5 5.5 30.5 6.5 ;
      RECT 29.5 31.5 30.5 32.5 ;
      RECT 29.5 33.5 30.5 34.5 ;
      RECT 25.5 5.5 26.5 6.5 ;
      RECT 25.5 13.5 26.5 14.5 ;
      RECT 25.5 31.5 26.5 32.5 ;
      RECT 25.5 33.5 26.5 34.5 ;
      RECT 21.5 5.5 22.5 6.5 ;
      RECT 21.5 31.5 22.5 32.5 ;
      RECT 21.5 33.5 22.5 34.5 ;
      RECT 17.5 5.5 18.5 6.5 ;
      RECT 17.5 17.5 18.5 18.5 ;
      RECT 17.5 31.5 18.5 32.5 ;
      RECT 17.5 33.5 18.5 34.5 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 17.5 14.5 18.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 25.5 2.5 26.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END AND4X1

MACRO AO21X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21X1 0 0 ;
  SIZE 32 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 32 3 ;
        RECT 25 -3 27 7 ;
        RECT 21 -3 23 7 ;
        RECT 1 -3 3 7 ;
    END
  END VSS!
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 13 9 15 15 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 29 5 31 31 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 17 9 19 15 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 13 3 19 ;
    END
  END C
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 32 43 ;
        RECT 25 27 27 43 ;
        RECT 1 27 3 43 ;
    END
  END VDD!
  PIN YN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9 17 27 19 ;
        RECT 21 17 23 31 ;
        RECT 9 5 11 31 ;
        RECT 5 5 11 7 ;
    END
  END YN
  OBS
    LAYER Metal1 ;
      RECT 5 33 19 35 ;
      RECT 17 27 19 35 ;
      RECT 13 27 15 35 ;
      RECT 5 27 7 35 ;
      RECT 13 5 19 7 ;
    LAYER Via1 ;
      RECT 29.5 5.5 30.5 6.5 ;
      RECT 29.5 27.5 30.5 28.5 ;
      RECT 29.5 29.5 30.5 30.5 ;
      RECT 25.5 5.5 26.5 6.5 ;
      RECT 25.5 17.5 26.5 18.5 ;
      RECT 25.5 27.5 26.5 28.5 ;
      RECT 25.5 29.5 26.5 30.5 ;
      RECT 21.5 5.5 22.5 6.5 ;
      RECT 21.5 27.5 22.5 28.5 ;
      RECT 21.5 29.5 22.5 30.5 ;
      RECT 17.5 5.5 18.5 6.5 ;
      RECT 17.5 13.5 18.5 14.5 ;
      RECT 17.5 27.5 18.5 28.5 ;
      RECT 17.5 29.5 18.5 30.5 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 9.5 14.5 10.5 ;
      RECT 13.5 27.5 14.5 28.5 ;
      RECT 13.5 29.5 14.5 30.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 27.5 10.5 28.5 ;
      RECT 9.5 29.5 10.5 30.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 27.5 6.5 28.5 ;
      RECT 5.5 29.5 6.5 30.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 13.5 2.5 14.5 ;
      RECT 1.5 27.5 2.5 28.5 ;
      RECT 1.5 29.5 2.5 30.5 ;
  END
END AO21X1

MACRO AOI21X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21X1 0 0 ;
  SIZE 24 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 24 3 ;
        RECT 21 -3 23 7 ;
        RECT 1 -3 3 7 ;
    END
  END VSS!
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 13 9 15 15 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 21 17 23 31 ;
        RECT 9 17 23 19 ;
        RECT 9 5 11 31 ;
        RECT 5 5 11 7 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 17 9 19 15 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 13 3 19 ;
    END
  END C
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 24 43 ;
        RECT 1 27 3 43 ;
    END
  END VDD!
  OBS
    LAYER Metal1 ;
      RECT 5 33 19 35 ;
      RECT 17 27 19 35 ;
      RECT 13 27 15 35 ;
      RECT 5 27 7 35 ;
      RECT 13 5 19 7 ;
    LAYER Via1 ;
      RECT 21.5 5.5 22.5 6.5 ;
      RECT 21.5 27.5 22.5 28.5 ;
      RECT 21.5 29.5 22.5 30.5 ;
      RECT 17.5 5.5 18.5 6.5 ;
      RECT 17.5 13.5 18.5 14.5 ;
      RECT 17.5 27.5 18.5 28.5 ;
      RECT 17.5 29.5 18.5 30.5 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 9.5 14.5 10.5 ;
      RECT 13.5 27.5 14.5 28.5 ;
      RECT 13.5 29.5 14.5 30.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 27.5 10.5 28.5 ;
      RECT 9.5 29.5 10.5 30.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 27.5 6.5 28.5 ;
      RECT 5.5 29.5 6.5 30.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 13.5 2.5 14.5 ;
      RECT 1.5 27.5 2.5 28.5 ;
      RECT 1.5 29.5 2.5 30.5 ;
  END
END AOI21X1

MACRO BUFX16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX16 0 0 ;
  SIZE 56 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 56 43 ;
        RECT 53 27 55 43 ;
        RECT 45 27 47 43 ;
        RECT 37 27 39 43 ;
        RECT 29 27 31 43 ;
        RECT 21 27 23 43 ;
        RECT 17 27 19 43 ;
        RECT 9 27 11 43 ;
        RECT 1 27 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 13 3 19 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 49 5 51 35 ;
        RECT 25 17 51 19 ;
        RECT 41 5 43 35 ;
        RECT 33 5 35 35 ;
        RECT 25 5 27 35 ;
    END
  END Y
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 56 3 ;
        RECT 53 -3 55 9 ;
        RECT 45 -3 47 9 ;
        RECT 37 -3 39 9 ;
        RECT 29 -3 31 9 ;
        RECT 21 -3 23 9 ;
        RECT 17 -3 19 9 ;
        RECT 9 -3 11 9 ;
        RECT 1 -3 3 9 ;
    END
  END VSS!
  OBS
    LAYER Metal1 ;
      RECT 13 5 15 35 ;
      RECT 5 5 7 35 ;
      RECT 5 13 23 15 ;
    LAYER Via1 ;
      RECT 53.5 5.5 54.5 6.5 ;
      RECT 53.5 7.5 54.5 8.5 ;
      RECT 53.5 27.5 54.5 28.5 ;
      RECT 53.5 29.5 54.5 30.5 ;
      RECT 53.5 31.5 54.5 32.5 ;
      RECT 53.5 33.5 54.5 34.5 ;
      RECT 49.5 5.5 50.5 6.5 ;
      RECT 49.5 7.5 50.5 8.5 ;
      RECT 49.5 27.5 50.5 28.5 ;
      RECT 49.5 29.5 50.5 30.5 ;
      RECT 49.5 31.5 50.5 32.5 ;
      RECT 49.5 33.5 50.5 34.5 ;
      RECT 45.5 5.5 46.5 6.5 ;
      RECT 45.5 7.5 46.5 8.5 ;
      RECT 45.5 27.5 46.5 28.5 ;
      RECT 45.5 29.5 46.5 30.5 ;
      RECT 45.5 31.5 46.5 32.5 ;
      RECT 45.5 33.5 46.5 34.5 ;
      RECT 41.5 5.5 42.5 6.5 ;
      RECT 41.5 7.5 42.5 8.5 ;
      RECT 41.5 27.5 42.5 28.5 ;
      RECT 41.5 29.5 42.5 30.5 ;
      RECT 41.5 31.5 42.5 32.5 ;
      RECT 41.5 33.5 42.5 34.5 ;
      RECT 37.5 5.5 38.5 6.5 ;
      RECT 37.5 7.5 38.5 8.5 ;
      RECT 37.5 27.5 38.5 28.5 ;
      RECT 37.5 29.5 38.5 30.5 ;
      RECT 37.5 31.5 38.5 32.5 ;
      RECT 37.5 33.5 38.5 34.5 ;
      RECT 33.5 5.5 34.5 6.5 ;
      RECT 33.5 7.5 34.5 8.5 ;
      RECT 33.5 27.5 34.5 28.5 ;
      RECT 33.5 29.5 34.5 30.5 ;
      RECT 33.5 31.5 34.5 32.5 ;
      RECT 33.5 33.5 34.5 34.5 ;
      RECT 29.5 5.5 30.5 6.5 ;
      RECT 29.5 7.5 30.5 8.5 ;
      RECT 29.5 27.5 30.5 28.5 ;
      RECT 29.5 29.5 30.5 30.5 ;
      RECT 29.5 31.5 30.5 32.5 ;
      RECT 29.5 33.5 30.5 34.5 ;
      RECT 25.5 5.5 26.5 6.5 ;
      RECT 25.5 7.5 26.5 8.5 ;
      RECT 25.5 27.5 26.5 28.5 ;
      RECT 25.5 29.5 26.5 30.5 ;
      RECT 25.5 31.5 26.5 32.5 ;
      RECT 25.5 33.5 26.5 34.5 ;
      RECT 21.5 5.5 22.5 6.5 ;
      RECT 21.5 7.5 22.5 8.5 ;
      RECT 21.5 13.5 22.5 14.5 ;
      RECT 21.5 27.5 22.5 28.5 ;
      RECT 21.5 29.5 22.5 30.5 ;
      RECT 21.5 31.5 22.5 32.5 ;
      RECT 21.5 33.5 22.5 34.5 ;
      RECT 17.5 5.5 18.5 6.5 ;
      RECT 17.5 7.5 18.5 8.5 ;
      RECT 17.5 27.5 18.5 28.5 ;
      RECT 17.5 29.5 18.5 30.5 ;
      RECT 17.5 31.5 18.5 32.5 ;
      RECT 17.5 33.5 18.5 34.5 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 7.5 14.5 8.5 ;
      RECT 13.5 27.5 14.5 28.5 ;
      RECT 13.5 29.5 14.5 30.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 7.5 10.5 8.5 ;
      RECT 9.5 27.5 10.5 28.5 ;
      RECT 9.5 29.5 10.5 30.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 7.5 6.5 8.5 ;
      RECT 5.5 27.5 6.5 28.5 ;
      RECT 5.5 29.5 6.5 30.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 7.5 2.5 8.5 ;
      RECT 1.5 17.5 2.5 18.5 ;
      RECT 1.5 27.5 2.5 28.5 ;
      RECT 1.5 29.5 2.5 30.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END BUFX16

MACRO BUFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX2 0 0 ;
  SIZE 16 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 16 43 ;
        RECT 9 27 11 43 ;
        RECT 1 31 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 17 3 23 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 13 5 15 35 ;
    END
  END Y
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 16 3 ;
        RECT 9 -3 11 9 ;
        RECT 1 -3 3 7 ;
    END
  END VSS!
  OBS
    LAYER Metal1 ;
      RECT 5 5 7 35 ;
      RECT 5 17 11 19 ;
    LAYER Via1 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 7.5 14.5 8.5 ;
      RECT 13.5 27.5 14.5 28.5 ;
      RECT 13.5 29.5 14.5 30.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 7.5 10.5 8.5 ;
      RECT 9.5 17.5 10.5 18.5 ;
      RECT 9.5 27.5 10.5 28.5 ;
      RECT 9.5 29.5 10.5 30.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 21.5 2.5 22.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END BUFX2

MACRO BUFX27
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX27 0 0 ;
  SIZE 56 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 56 43 ;
        RECT 49 23 51 43 ;
        RECT 41 23 43 43 ;
        RECT 33 23 35 43 ;
        RECT 25 23 27 43 ;
        RECT 17 23 19 43 ;
        RECT 9 23 11 43 ;
        RECT 1 23 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 13 3 19 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 53 5 55 35 ;
        RECT 21 13 55 15 ;
        RECT 45 5 47 35 ;
        RECT 37 5 39 35 ;
        RECT 29 5 31 35 ;
        RECT 21 5 23 35 ;
    END
  END Y
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 56 3 ;
        RECT 49 -3 51 11 ;
        RECT 41 -3 43 11 ;
        RECT 33 -3 35 11 ;
        RECT 25 -3 27 11 ;
        RECT 17 -3 19 11 ;
        RECT 9 -3 11 11 ;
        RECT 1 -3 3 11 ;
    END
  END VSS!
  OBS
    LAYER Metal1 ;
      RECT 13 5 15 35 ;
      RECT 5 5 7 35 ;
      RECT 5 17 19 19 ;
    LAYER Via1 ;
      RECT 53.5 5.5 54.5 6.5 ;
      RECT 53.5 7.5 54.5 8.5 ;
      RECT 53.5 9.5 54.5 10.5 ;
      RECT 53.5 23.5 54.5 24.5 ;
      RECT 53.5 25.5 54.5 26.5 ;
      RECT 53.5 27.5 54.5 28.5 ;
      RECT 53.5 29.5 54.5 30.5 ;
      RECT 53.5 31.5 54.5 32.5 ;
      RECT 53.5 33.5 54.5 34.5 ;
      RECT 49.5 5.5 50.5 6.5 ;
      RECT 49.5 7.5 50.5 8.5 ;
      RECT 49.5 9.5 50.5 10.5 ;
      RECT 49.5 23.5 50.5 24.5 ;
      RECT 49.5 25.5 50.5 26.5 ;
      RECT 49.5 27.5 50.5 28.5 ;
      RECT 49.5 29.5 50.5 30.5 ;
      RECT 49.5 31.5 50.5 32.5 ;
      RECT 49.5 33.5 50.5 34.5 ;
      RECT 45.5 5.5 46.5 6.5 ;
      RECT 45.5 7.5 46.5 8.5 ;
      RECT 45.5 9.5 46.5 10.5 ;
      RECT 45.5 23.5 46.5 24.5 ;
      RECT 45.5 25.5 46.5 26.5 ;
      RECT 45.5 27.5 46.5 28.5 ;
      RECT 45.5 29.5 46.5 30.5 ;
      RECT 45.5 31.5 46.5 32.5 ;
      RECT 45.5 33.5 46.5 34.5 ;
      RECT 41.5 5.5 42.5 6.5 ;
      RECT 41.5 7.5 42.5 8.5 ;
      RECT 41.5 9.5 42.5 10.5 ;
      RECT 41.5 23.5 42.5 24.5 ;
      RECT 41.5 25.5 42.5 26.5 ;
      RECT 41.5 27.5 42.5 28.5 ;
      RECT 41.5 29.5 42.5 30.5 ;
      RECT 41.5 31.5 42.5 32.5 ;
      RECT 41.5 33.5 42.5 34.5 ;
      RECT 37.5 5.5 38.5 6.5 ;
      RECT 37.5 7.5 38.5 8.5 ;
      RECT 37.5 9.5 38.5 10.5 ;
      RECT 37.5 23.5 38.5 24.5 ;
      RECT 37.5 25.5 38.5 26.5 ;
      RECT 37.5 27.5 38.5 28.5 ;
      RECT 37.5 29.5 38.5 30.5 ;
      RECT 37.5 31.5 38.5 32.5 ;
      RECT 37.5 33.5 38.5 34.5 ;
      RECT 33.5 5.5 34.5 6.5 ;
      RECT 33.5 7.5 34.5 8.5 ;
      RECT 33.5 9.5 34.5 10.5 ;
      RECT 33.5 23.5 34.5 24.5 ;
      RECT 33.5 25.5 34.5 26.5 ;
      RECT 33.5 27.5 34.5 28.5 ;
      RECT 33.5 29.5 34.5 30.5 ;
      RECT 33.5 31.5 34.5 32.5 ;
      RECT 33.5 33.5 34.5 34.5 ;
      RECT 29.5 5.5 30.5 6.5 ;
      RECT 29.5 7.5 30.5 8.5 ;
      RECT 29.5 9.5 30.5 10.5 ;
      RECT 29.5 23.5 30.5 24.5 ;
      RECT 29.5 25.5 30.5 26.5 ;
      RECT 29.5 27.5 30.5 28.5 ;
      RECT 29.5 29.5 30.5 30.5 ;
      RECT 29.5 31.5 30.5 32.5 ;
      RECT 29.5 33.5 30.5 34.5 ;
      RECT 25.5 5.5 26.5 6.5 ;
      RECT 25.5 7.5 26.5 8.5 ;
      RECT 25.5 9.5 26.5 10.5 ;
      RECT 25.5 23.5 26.5 24.5 ;
      RECT 25.5 25.5 26.5 26.5 ;
      RECT 25.5 27.5 26.5 28.5 ;
      RECT 25.5 29.5 26.5 30.5 ;
      RECT 25.5 31.5 26.5 32.5 ;
      RECT 25.5 33.5 26.5 34.5 ;
      RECT 21.5 5.5 22.5 6.5 ;
      RECT 21.5 7.5 22.5 8.5 ;
      RECT 21.5 9.5 22.5 10.5 ;
      RECT 21.5 23.5 22.5 24.5 ;
      RECT 21.5 25.5 22.5 26.5 ;
      RECT 21.5 27.5 22.5 28.5 ;
      RECT 21.5 29.5 22.5 30.5 ;
      RECT 21.5 31.5 22.5 32.5 ;
      RECT 21.5 33.5 22.5 34.5 ;
      RECT 17.5 5.5 18.5 6.5 ;
      RECT 17.5 7.5 18.5 8.5 ;
      RECT 17.5 9.5 18.5 10.5 ;
      RECT 17.5 17.5 18.5 18.5 ;
      RECT 17.5 23.5 18.5 24.5 ;
      RECT 17.5 25.5 18.5 26.5 ;
      RECT 17.5 27.5 18.5 28.5 ;
      RECT 17.5 29.5 18.5 30.5 ;
      RECT 17.5 31.5 18.5 32.5 ;
      RECT 17.5 33.5 18.5 34.5 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 7.5 14.5 8.5 ;
      RECT 13.5 9.5 14.5 10.5 ;
      RECT 13.5 23.5 14.5 24.5 ;
      RECT 13.5 25.5 14.5 26.5 ;
      RECT 13.5 27.5 14.5 28.5 ;
      RECT 13.5 29.5 14.5 30.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 7.5 10.5 8.5 ;
      RECT 9.5 9.5 10.5 10.5 ;
      RECT 9.5 23.5 10.5 24.5 ;
      RECT 9.5 25.5 10.5 26.5 ;
      RECT 9.5 27.5 10.5 28.5 ;
      RECT 9.5 29.5 10.5 30.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 7.5 6.5 8.5 ;
      RECT 5.5 9.5 6.5 10.5 ;
      RECT 5.5 23.5 6.5 24.5 ;
      RECT 5.5 25.5 6.5 26.5 ;
      RECT 5.5 27.5 6.5 28.5 ;
      RECT 5.5 29.5 6.5 30.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 7.5 2.5 8.5 ;
      RECT 1.5 9.5 2.5 10.5 ;
      RECT 1.5 13.5 2.5 14.5 ;
      RECT 1.5 23.5 2.5 24.5 ;
      RECT 1.5 25.5 2.5 26.5 ;
      RECT 1.5 27.5 2.5 28.5 ;
      RECT 1.5 29.5 2.5 30.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END BUFX27

MACRO BUFX3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX3 0 0 ;
  SIZE 16 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 16 43 ;
        RECT 9 23 11 43 ;
        RECT 1 31 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 21 3 27 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 13 5 15 35 ;
    END
  END Y
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 16 3 ;
        RECT 9 -3 11 11 ;
        RECT 1 -3 3 7 ;
    END
  END VSS!
  OBS
    LAYER Metal1 ;
      RECT 5 5 7 35 ;
      RECT 5 13 11 15 ;
    LAYER Via1 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 7.5 14.5 8.5 ;
      RECT 13.5 9.5 14.5 10.5 ;
      RECT 13.5 23.5 14.5 24.5 ;
      RECT 13.5 25.5 14.5 26.5 ;
      RECT 13.5 27.5 14.5 28.5 ;
      RECT 13.5 29.5 14.5 30.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 7.5 10.5 8.5 ;
      RECT 9.5 9.5 10.5 10.5 ;
      RECT 9.5 13.5 10.5 14.5 ;
      RECT 9.5 23.5 10.5 24.5 ;
      RECT 9.5 25.5 10.5 26.5 ;
      RECT 9.5 27.5 10.5 28.5 ;
      RECT 9.5 29.5 10.5 30.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 25.5 2.5 26.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END BUFX3

MACRO BUFX32
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX32 0 0 ;
  SIZE 104 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 104 43 ;
        RECT 101 27 103 43 ;
        RECT 93 27 95 43 ;
        RECT 85 27 87 43 ;
        RECT 77 27 79 43 ;
        RECT 69 27 71 43 ;
        RECT 61 27 63 43 ;
        RECT 53 27 55 43 ;
        RECT 45 27 47 43 ;
        RECT 37 27 39 43 ;
        RECT 33 27 35 43 ;
        RECT 25 27 27 43 ;
        RECT 17 27 19 43 ;
        RECT 9 27 11 43 ;
        RECT 1 27 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 13 3 19 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 97 5 99 35 ;
        RECT 41 17 99 19 ;
        RECT 89 5 91 35 ;
        RECT 81 5 83 35 ;
        RECT 73 5 75 35 ;
        RECT 65 5 67 35 ;
        RECT 57 5 59 35 ;
        RECT 49 5 51 35 ;
        RECT 41 5 43 35 ;
    END
  END Y
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 104 3 ;
        RECT 101 -3 103 9 ;
        RECT 93 -3 95 9 ;
        RECT 85 -3 87 9 ;
        RECT 77 -3 79 9 ;
        RECT 69 -3 71 9 ;
        RECT 61 -3 63 9 ;
        RECT 53 -3 55 9 ;
        RECT 45 -3 47 9 ;
        RECT 37 -3 39 9 ;
        RECT 33 -3 35 9 ;
        RECT 25 -3 27 9 ;
        RECT 17 -3 19 9 ;
        RECT 9 -3 11 9 ;
        RECT 1 -3 3 9 ;
    END
  END VSS!
  OBS
    LAYER Metal1 ;
      RECT 29 5 31 35 ;
      RECT 21 5 23 35 ;
      RECT 13 5 15 35 ;
      RECT 5 5 7 35 ;
      RECT 5 13 39 15 ;
    LAYER Via1 ;
      RECT 101.5 5.5 102.5 6.5 ;
      RECT 101.5 7.5 102.5 8.5 ;
      RECT 101.5 27.5 102.5 28.5 ;
      RECT 101.5 29.5 102.5 30.5 ;
      RECT 101.5 31.5 102.5 32.5 ;
      RECT 101.5 33.5 102.5 34.5 ;
      RECT 97.5 5.5 98.5 6.5 ;
      RECT 97.5 7.5 98.5 8.5 ;
      RECT 97.5 27.5 98.5 28.5 ;
      RECT 97.5 29.5 98.5 30.5 ;
      RECT 97.5 31.5 98.5 32.5 ;
      RECT 97.5 33.5 98.5 34.5 ;
      RECT 93.5 5.5 94.5 6.5 ;
      RECT 93.5 7.5 94.5 8.5 ;
      RECT 93.5 27.5 94.5 28.5 ;
      RECT 93.5 29.5 94.5 30.5 ;
      RECT 93.5 31.5 94.5 32.5 ;
      RECT 93.5 33.5 94.5 34.5 ;
      RECT 89.5 5.5 90.5 6.5 ;
      RECT 89.5 7.5 90.5 8.5 ;
      RECT 89.5 27.5 90.5 28.5 ;
      RECT 89.5 29.5 90.5 30.5 ;
      RECT 89.5 31.5 90.5 32.5 ;
      RECT 89.5 33.5 90.5 34.5 ;
      RECT 85.5 5.5 86.5 6.5 ;
      RECT 85.5 7.5 86.5 8.5 ;
      RECT 85.5 27.5 86.5 28.5 ;
      RECT 85.5 29.5 86.5 30.5 ;
      RECT 85.5 31.5 86.5 32.5 ;
      RECT 85.5 33.5 86.5 34.5 ;
      RECT 81.5 5.5 82.5 6.5 ;
      RECT 81.5 7.5 82.5 8.5 ;
      RECT 81.5 27.5 82.5 28.5 ;
      RECT 81.5 29.5 82.5 30.5 ;
      RECT 81.5 31.5 82.5 32.5 ;
      RECT 81.5 33.5 82.5 34.5 ;
      RECT 77.5 5.5 78.5 6.5 ;
      RECT 77.5 7.5 78.5 8.5 ;
      RECT 77.5 27.5 78.5 28.5 ;
      RECT 77.5 29.5 78.5 30.5 ;
      RECT 77.5 31.5 78.5 32.5 ;
      RECT 77.5 33.5 78.5 34.5 ;
      RECT 73.5 5.5 74.5 6.5 ;
      RECT 73.5 7.5 74.5 8.5 ;
      RECT 73.5 27.5 74.5 28.5 ;
      RECT 73.5 29.5 74.5 30.5 ;
      RECT 73.5 31.5 74.5 32.5 ;
      RECT 73.5 33.5 74.5 34.5 ;
      RECT 69.5 5.5 70.5 6.5 ;
      RECT 69.5 7.5 70.5 8.5 ;
      RECT 69.5 27.5 70.5 28.5 ;
      RECT 69.5 29.5 70.5 30.5 ;
      RECT 69.5 31.5 70.5 32.5 ;
      RECT 69.5 33.5 70.5 34.5 ;
      RECT 65.5 5.5 66.5 6.5 ;
      RECT 65.5 7.5 66.5 8.5 ;
      RECT 65.5 27.5 66.5 28.5 ;
      RECT 65.5 29.5 66.5 30.5 ;
      RECT 65.5 31.5 66.5 32.5 ;
      RECT 65.5 33.5 66.5 34.5 ;
      RECT 61.5 5.5 62.5 6.5 ;
      RECT 61.5 7.5 62.5 8.5 ;
      RECT 61.5 27.5 62.5 28.5 ;
      RECT 61.5 29.5 62.5 30.5 ;
      RECT 61.5 31.5 62.5 32.5 ;
      RECT 61.5 33.5 62.5 34.5 ;
      RECT 57.5 5.5 58.5 6.5 ;
      RECT 57.5 7.5 58.5 8.5 ;
      RECT 57.5 27.5 58.5 28.5 ;
      RECT 57.5 29.5 58.5 30.5 ;
      RECT 57.5 31.5 58.5 32.5 ;
      RECT 57.5 33.5 58.5 34.5 ;
      RECT 53.5 5.5 54.5 6.5 ;
      RECT 53.5 7.5 54.5 8.5 ;
      RECT 53.5 27.5 54.5 28.5 ;
      RECT 53.5 29.5 54.5 30.5 ;
      RECT 53.5 31.5 54.5 32.5 ;
      RECT 53.5 33.5 54.5 34.5 ;
      RECT 49.5 5.5 50.5 6.5 ;
      RECT 49.5 7.5 50.5 8.5 ;
      RECT 49.5 27.5 50.5 28.5 ;
      RECT 49.5 29.5 50.5 30.5 ;
      RECT 49.5 31.5 50.5 32.5 ;
      RECT 49.5 33.5 50.5 34.5 ;
      RECT 45.5 5.5 46.5 6.5 ;
      RECT 45.5 7.5 46.5 8.5 ;
      RECT 45.5 27.5 46.5 28.5 ;
      RECT 45.5 29.5 46.5 30.5 ;
      RECT 45.5 31.5 46.5 32.5 ;
      RECT 45.5 33.5 46.5 34.5 ;
      RECT 41.5 5.5 42.5 6.5 ;
      RECT 41.5 7.5 42.5 8.5 ;
      RECT 41.5 27.5 42.5 28.5 ;
      RECT 41.5 29.5 42.5 30.5 ;
      RECT 41.5 31.5 42.5 32.5 ;
      RECT 41.5 33.5 42.5 34.5 ;
      RECT 37.5 5.5 38.5 6.5 ;
      RECT 37.5 7.5 38.5 8.5 ;
      RECT 37.5 13.5 38.5 14.5 ;
      RECT 37.5 27.5 38.5 28.5 ;
      RECT 37.5 29.5 38.5 30.5 ;
      RECT 37.5 31.5 38.5 32.5 ;
      RECT 37.5 33.5 38.5 34.5 ;
      RECT 33.5 5.5 34.5 6.5 ;
      RECT 33.5 7.5 34.5 8.5 ;
      RECT 33.5 27.5 34.5 28.5 ;
      RECT 33.5 29.5 34.5 30.5 ;
      RECT 33.5 31.5 34.5 32.5 ;
      RECT 33.5 33.5 34.5 34.5 ;
      RECT 29.5 5.5 30.5 6.5 ;
      RECT 29.5 7.5 30.5 8.5 ;
      RECT 29.5 27.5 30.5 28.5 ;
      RECT 29.5 29.5 30.5 30.5 ;
      RECT 29.5 31.5 30.5 32.5 ;
      RECT 29.5 33.5 30.5 34.5 ;
      RECT 25.5 5.5 26.5 6.5 ;
      RECT 25.5 7.5 26.5 8.5 ;
      RECT 25.5 27.5 26.5 28.5 ;
      RECT 25.5 29.5 26.5 30.5 ;
      RECT 25.5 31.5 26.5 32.5 ;
      RECT 25.5 33.5 26.5 34.5 ;
      RECT 21.5 5.5 22.5 6.5 ;
      RECT 21.5 7.5 22.5 8.5 ;
      RECT 21.5 27.5 22.5 28.5 ;
      RECT 21.5 29.5 22.5 30.5 ;
      RECT 21.5 31.5 22.5 32.5 ;
      RECT 21.5 33.5 22.5 34.5 ;
      RECT 17.5 5.5 18.5 6.5 ;
      RECT 17.5 7.5 18.5 8.5 ;
      RECT 17.5 27.5 18.5 28.5 ;
      RECT 17.5 29.5 18.5 30.5 ;
      RECT 17.5 31.5 18.5 32.5 ;
      RECT 17.5 33.5 18.5 34.5 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 7.5 14.5 8.5 ;
      RECT 13.5 27.5 14.5 28.5 ;
      RECT 13.5 29.5 14.5 30.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 7.5 10.5 8.5 ;
      RECT 9.5 27.5 10.5 28.5 ;
      RECT 9.5 29.5 10.5 30.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 7.5 6.5 8.5 ;
      RECT 5.5 27.5 6.5 28.5 ;
      RECT 5.5 29.5 6.5 30.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 7.5 2.5 8.5 ;
      RECT 1.5 17.5 2.5 18.5 ;
      RECT 1.5 27.5 2.5 28.5 ;
      RECT 1.5 29.5 2.5 30.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END BUFX32

MACRO BUFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX4 0 0 ;
  SIZE 20 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 20 43 ;
        RECT 17 27 19 43 ;
        RECT 9 27 11 43 ;
        RECT 1 27 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 13 3 19 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 13 5 15 35 ;
    END
  END Y
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 20 3 ;
        RECT 17 -3 19 9 ;
        RECT 9 -3 11 9 ;
        RECT 1 -3 3 9 ;
    END
  END VSS!
  OBS
    LAYER Metal1 ;
      RECT 5 5 7 35 ;
      RECT 5 17 11 19 ;
    LAYER Via1 ;
      RECT 17.5 5.5 18.5 6.5 ;
      RECT 17.5 7.5 18.5 8.5 ;
      RECT 17.5 27.5 18.5 28.5 ;
      RECT 17.5 29.5 18.5 30.5 ;
      RECT 17.5 31.5 18.5 32.5 ;
      RECT 17.5 33.5 18.5 34.5 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 7.5 14.5 8.5 ;
      RECT 13.5 27.5 14.5 28.5 ;
      RECT 13.5 29.5 14.5 30.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 7.5 10.5 8.5 ;
      RECT 9.5 17.5 10.5 18.5 ;
      RECT 9.5 27.5 10.5 28.5 ;
      RECT 9.5 29.5 10.5 30.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 7.5 6.5 8.5 ;
      RECT 5.5 27.5 6.5 28.5 ;
      RECT 5.5 29.5 6.5 30.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 7.5 2.5 8.5 ;
      RECT 1.5 17.5 2.5 18.5 ;
      RECT 1.5 27.5 2.5 28.5 ;
      RECT 1.5 29.5 2.5 30.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END BUFX4

MACRO BUFX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX8 0 0 ;
  SIZE 32 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 32 43 ;
        RECT 29 27 31 43 ;
        RECT 21 27 23 43 ;
        RECT 13 27 15 43 ;
        RECT 9 27 11 43 ;
        RECT 1 27 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 13 3 19 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 25 5 27 35 ;
        RECT 17 17 27 19 ;
        RECT 17 5 19 35 ;
    END
  END Y
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 32 3 ;
        RECT 29 -3 31 9 ;
        RECT 21 -3 23 9 ;
        RECT 13 -3 15 9 ;
        RECT 9 -3 11 9 ;
        RECT 1 -3 3 9 ;
    END
  END VSS!
  OBS
    LAYER Metal1 ;
      RECT 5 5 7 35 ;
      RECT 5 13 15 15 ;
    LAYER Via1 ;
      RECT 29.5 5.5 30.5 6.5 ;
      RECT 29.5 7.5 30.5 8.5 ;
      RECT 29.5 27.5 30.5 28.5 ;
      RECT 29.5 29.5 30.5 30.5 ;
      RECT 29.5 31.5 30.5 32.5 ;
      RECT 29.5 33.5 30.5 34.5 ;
      RECT 25.5 5.5 26.5 6.5 ;
      RECT 25.5 7.5 26.5 8.5 ;
      RECT 25.5 27.5 26.5 28.5 ;
      RECT 25.5 29.5 26.5 30.5 ;
      RECT 25.5 31.5 26.5 32.5 ;
      RECT 25.5 33.5 26.5 34.5 ;
      RECT 21.5 5.5 22.5 6.5 ;
      RECT 21.5 7.5 22.5 8.5 ;
      RECT 21.5 27.5 22.5 28.5 ;
      RECT 21.5 29.5 22.5 30.5 ;
      RECT 21.5 31.5 22.5 32.5 ;
      RECT 21.5 33.5 22.5 34.5 ;
      RECT 17.5 5.5 18.5 6.5 ;
      RECT 17.5 7.5 18.5 8.5 ;
      RECT 17.5 27.5 18.5 28.5 ;
      RECT 17.5 29.5 18.5 30.5 ;
      RECT 17.5 31.5 18.5 32.5 ;
      RECT 17.5 33.5 18.5 34.5 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 7.5 14.5 8.5 ;
      RECT 13.5 13.5 14.5 14.5 ;
      RECT 13.5 27.5 14.5 28.5 ;
      RECT 13.5 29.5 14.5 30.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 7.5 10.5 8.5 ;
      RECT 9.5 27.5 10.5 28.5 ;
      RECT 9.5 29.5 10.5 30.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 7.5 6.5 8.5 ;
      RECT 5.5 27.5 6.5 28.5 ;
      RECT 5.5 29.5 6.5 30.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 7.5 2.5 8.5 ;
      RECT 1.5 17.5 2.5 18.5 ;
      RECT 1.5 27.5 2.5 28.5 ;
      RECT 1.5 29.5 2.5 30.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END BUFX8

MACRO BUFX9
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX9 0 0 ;
  SIZE 24 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 24 43 ;
        RECT 17 23 19 43 ;
        RECT 9 23 11 43 ;
        RECT 1 23 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 13 3 19 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 21 5 23 35 ;
        RECT 13 17 23 19 ;
        RECT 13 5 15 35 ;
    END
  END Y
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 24 3 ;
        RECT 17 -3 19 11 ;
        RECT 9 -3 11 11 ;
        RECT 1 -3 3 11 ;
    END
  END VSS!
  OBS
    LAYER Metal1 ;
      RECT 5 5 7 35 ;
      RECT 5 13 11 15 ;
    LAYER Via1 ;
      RECT 21.5 5.5 22.5 6.5 ;
      RECT 21.5 7.5 22.5 8.5 ;
      RECT 21.5 9.5 22.5 10.5 ;
      RECT 21.5 23.5 22.5 24.5 ;
      RECT 21.5 25.5 22.5 26.5 ;
      RECT 21.5 27.5 22.5 28.5 ;
      RECT 21.5 29.5 22.5 30.5 ;
      RECT 21.5 31.5 22.5 32.5 ;
      RECT 21.5 33.5 22.5 34.5 ;
      RECT 17.5 5.5 18.5 6.5 ;
      RECT 17.5 7.5 18.5 8.5 ;
      RECT 17.5 9.5 18.5 10.5 ;
      RECT 17.5 23.5 18.5 24.5 ;
      RECT 17.5 25.5 18.5 26.5 ;
      RECT 17.5 27.5 18.5 28.5 ;
      RECT 17.5 29.5 18.5 30.5 ;
      RECT 17.5 31.5 18.5 32.5 ;
      RECT 17.5 33.5 18.5 34.5 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 7.5 14.5 8.5 ;
      RECT 13.5 9.5 14.5 10.5 ;
      RECT 13.5 23.5 14.5 24.5 ;
      RECT 13.5 25.5 14.5 26.5 ;
      RECT 13.5 27.5 14.5 28.5 ;
      RECT 13.5 29.5 14.5 30.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 7.5 10.5 8.5 ;
      RECT 9.5 9.5 10.5 10.5 ;
      RECT 9.5 13.5 10.5 14.5 ;
      RECT 9.5 23.5 10.5 24.5 ;
      RECT 9.5 25.5 10.5 26.5 ;
      RECT 9.5 27.5 10.5 28.5 ;
      RECT 9.5 29.5 10.5 30.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 7.5 6.5 8.5 ;
      RECT 5.5 9.5 6.5 10.5 ;
      RECT 5.5 23.5 6.5 24.5 ;
      RECT 5.5 25.5 6.5 26.5 ;
      RECT 5.5 27.5 6.5 28.5 ;
      RECT 5.5 29.5 6.5 30.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 7.5 2.5 8.5 ;
      RECT 1.5 9.5 2.5 10.5 ;
      RECT 1.5 13.5 2.5 14.5 ;
      RECT 1.5 23.5 2.5 24.5 ;
      RECT 1.5 25.5 2.5 26.5 ;
      RECT 1.5 27.5 2.5 28.5 ;
      RECT 1.5 29.5 2.5 30.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END BUFX9

MACRO DECAP2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DECAP2 0 0 ;
  SIZE 8 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 8 43 ;
        RECT 1 25 3 43 ;
    END
  END VDD!
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 8 3 ;
        RECT 5 -3 7 15 ;
    END
  END VSS!
  OBS
    LAYER Metal1 ;
      RECT 5 17 7 35 ;
      RECT 1 5 3 23 ;
    LAYER Via1 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 7.5 6.5 8.5 ;
      RECT 5.5 9.5 6.5 10.5 ;
      RECT 5.5 11.5 6.5 12.5 ;
      RECT 5.5 13.5 6.5 14.5 ;
      RECT 5.5 17.5 6.5 18.5 ;
      RECT 5.5 25.5 6.5 26.5 ;
      RECT 5.5 27.5 6.5 28.5 ;
      RECT 5.5 29.5 6.5 30.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 7.5 2.5 8.5 ;
      RECT 1.5 9.5 2.5 10.5 ;
      RECT 1.5 11.5 2.5 12.5 ;
      RECT 1.5 13.5 2.5 14.5 ;
      RECT 1.5 21.5 2.5 22.5 ;
      RECT 1.5 25.5 2.5 26.5 ;
      RECT 1.5 27.5 2.5 28.5 ;
      RECT 1.5 29.5 2.5 30.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END DECAP2

MACRO DECAP3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DECAP3 0 0 ;
  SIZE 16 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 16 43 ;
        RECT 1 25 3 43 ;
    END
  END VDD!
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 16 3 ;
        RECT 13 -3 15 15 ;
    END
  END VSS!
  OBS
    LAYER Metal1 ;
      RECT 13 17 15 35 ;
      RECT 1 5 3 23 ;
    LAYER Via1 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 7.5 14.5 8.5 ;
      RECT 13.5 9.5 14.5 10.5 ;
      RECT 13.5 11.5 14.5 12.5 ;
      RECT 13.5 13.5 14.5 14.5 ;
      RECT 13.5 17.5 14.5 18.5 ;
      RECT 13.5 25.5 14.5 26.5 ;
      RECT 13.5 27.5 14.5 28.5 ;
      RECT 13.5 29.5 14.5 30.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 7.5 2.5 8.5 ;
      RECT 1.5 9.5 2.5 10.5 ;
      RECT 1.5 11.5 2.5 12.5 ;
      RECT 1.5 13.5 2.5 14.5 ;
      RECT 1.5 21.5 2.5 22.5 ;
      RECT 1.5 25.5 2.5 26.5 ;
      RECT 1.5 27.5 2.5 28.5 ;
      RECT 1.5 29.5 2.5 30.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END DECAP3

MACRO DECAP4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DECAP4 0 0 ;
  SIZE 32 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 32 43 ;
        RECT 1 25 3 43 ;
    END
  END VDD!
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 32 3 ;
        RECT 29 -3 31 15 ;
    END
  END VSS!
  OBS
    LAYER Metal1 ;
      RECT 29 17 31 35 ;
      RECT 1 5 3 23 ;
    LAYER Via1 ;
      RECT 29.5 5.5 30.5 6.5 ;
      RECT 29.5 7.5 30.5 8.5 ;
      RECT 29.5 9.5 30.5 10.5 ;
      RECT 29.5 11.5 30.5 12.5 ;
      RECT 29.5 13.5 30.5 14.5 ;
      RECT 29.5 17.5 30.5 18.5 ;
      RECT 29.5 25.5 30.5 26.5 ;
      RECT 29.5 27.5 30.5 28.5 ;
      RECT 29.5 29.5 30.5 30.5 ;
      RECT 29.5 31.5 30.5 32.5 ;
      RECT 29.5 33.5 30.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 7.5 2.5 8.5 ;
      RECT 1.5 9.5 2.5 10.5 ;
      RECT 1.5 11.5 2.5 12.5 ;
      RECT 1.5 13.5 2.5 14.5 ;
      RECT 1.5 21.5 2.5 22.5 ;
      RECT 1.5 25.5 2.5 26.5 ;
      RECT 1.5 27.5 2.5 28.5 ;
      RECT 1.5 29.5 2.5 30.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END DECAP4

MACRO DFFRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRX1 0 0 ;
  SIZE 136 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 136 43 ;
        RECT 129 31 131 43 ;
        RECT 121 31 123 43 ;
        RECT 113 31 115 43 ;
        RECT 109 31 111 43 ;
        RECT 101 31 103 43 ;
        RECT 93 31 95 43 ;
        RECT 85 31 87 43 ;
        RECT 73 31 75 43 ;
        RECT 65 31 67 43 ;
        RECT 53 31 55 43 ;
        RECT 45 31 47 43 ;
        RECT 33 31 35 43 ;
        RECT 25 31 27 43 ;
        RECT 17 31 19 43 ;
        RECT 13 31 15 43 ;
        RECT 5 31 7 43 ;
    END
  END VDD!
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 136 3 ;
        RECT 133 -3 135 19 ;
        RECT 89 -3 91 7 ;
        RECT 85 -3 87 7 ;
        RECT 41 -3 43 7 ;
        RECT 37 -3 39 7 ;
        RECT 1 -3 3 7 ;
    END
  END VSS!
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 29 9 99 11 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 125 5 127 11 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 41 25 59 27 ;
        RECT 49 25 51 35 ;
        RECT 41 25 43 35 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 77 31 83 35 ;
        RECT 77 25 79 35 ;
        RECT 61 25 79 27 ;
        RECT 69 25 71 35 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 37 13 131 15 ;
    END
  END RN
  OBS
    LAYER Metal1 ;
      RECT 133 21 135 35 ;
      RECT 125 21 127 35 ;
      RECT 117 21 119 35 ;
      RECT 5 21 135 23 ;
      RECT 113 17 115 23 ;
      RECT 105 25 107 35 ;
      RECT 97 25 99 35 ;
      RECT 89 25 91 35 ;
      RECT 85 25 115 27 ;
      RECT 37 25 39 35 ;
      RECT 29 25 31 35 ;
      RECT 21 25 23 35 ;
      RECT 13 25 39 27 ;
      RECT 21 5 23 11 ;
      RECT 21 5 27 7 ;
      RECT 17 5 19 11 ;
      RECT 13 5 19 7 ;
      RECT 9 25 11 35 ;
      RECT 1 13 3 35 ;
      RECT 1 25 11 27 ;
      RECT 1 13 19 15 ;
      RECT 13 9 15 15 ;
      RECT 9 5 11 11 ;
      RECT 5 5 11 7 ;
      RECT 125 17 131 19 ;
      RECT 117 17 123 19 ;
      RECT 109 5 115 7 ;
      RECT 101 5 107 7 ;
      RECT 93 5 99 7 ;
      RECT 13 17 91 19 ;
      RECT 77 5 83 7 ;
      RECT 69 5 75 7 ;
      RECT 61 5 67 7 ;
      RECT 53 5 59 7 ;
      RECT 45 5 51 7 ;
      RECT 29 5 35 7 ;
    LAYER Via1 ;
      RECT 133.5 17.5 134.5 18.5 ;
      RECT 133.5 31.5 134.5 32.5 ;
      RECT 133.5 33.5 134.5 34.5 ;
      RECT 129.5 13.5 130.5 14.5 ;
      RECT 129.5 17.5 130.5 18.5 ;
      RECT 129.5 31.5 130.5 32.5 ;
      RECT 129.5 33.5 130.5 34.5 ;
      RECT 125.5 9.5 126.5 10.5 ;
      RECT 125.5 17.5 126.5 18.5 ;
      RECT 125.5 31.5 126.5 32.5 ;
      RECT 125.5 33.5 126.5 34.5 ;
      RECT 121.5 17.5 122.5 18.5 ;
      RECT 121.5 31.5 122.5 32.5 ;
      RECT 121.5 33.5 122.5 34.5 ;
      RECT 117.5 17.5 118.5 18.5 ;
      RECT 117.5 31.5 118.5 32.5 ;
      RECT 117.5 33.5 118.5 34.5 ;
      RECT 113.5 5.5 114.5 6.5 ;
      RECT 113.5 17.5 114.5 18.5 ;
      RECT 113.5 25.5 114.5 26.5 ;
      RECT 113.5 31.5 114.5 32.5 ;
      RECT 113.5 33.5 114.5 34.5 ;
      RECT 109.5 5.5 110.5 6.5 ;
      RECT 109.5 31.5 110.5 32.5 ;
      RECT 109.5 33.5 110.5 34.5 ;
      RECT 105.5 5.5 106.5 6.5 ;
      RECT 105.5 21.5 106.5 22.5 ;
      RECT 105.5 31.5 106.5 32.5 ;
      RECT 105.5 33.5 106.5 34.5 ;
      RECT 101.5 5.5 102.5 6.5 ;
      RECT 101.5 31.5 102.5 32.5 ;
      RECT 101.5 33.5 102.5 34.5 ;
      RECT 97.5 5.5 98.5 6.5 ;
      RECT 97.5 9.5 98.5 10.5 ;
      RECT 97.5 31.5 98.5 32.5 ;
      RECT 97.5 33.5 98.5 34.5 ;
      RECT 93.5 5.5 94.5 6.5 ;
      RECT 93.5 31.5 94.5 32.5 ;
      RECT 93.5 33.5 94.5 34.5 ;
      RECT 89.5 5.5 90.5 6.5 ;
      RECT 89.5 17.5 90.5 18.5 ;
      RECT 89.5 31.5 90.5 32.5 ;
      RECT 89.5 33.5 90.5 34.5 ;
      RECT 85.5 5.5 86.5 6.5 ;
      RECT 85.5 25.5 86.5 26.5 ;
      RECT 85.5 31.5 86.5 32.5 ;
      RECT 85.5 33.5 86.5 34.5 ;
      RECT 81.5 5.5 82.5 6.5 ;
      RECT 81.5 31.5 82.5 32.5 ;
      RECT 81.5 33.5 82.5 34.5 ;
      RECT 77.5 5.5 78.5 6.5 ;
      RECT 77.5 13.5 78.5 14.5 ;
      RECT 77.5 31.5 78.5 32.5 ;
      RECT 77.5 33.5 78.5 34.5 ;
      RECT 73.5 5.5 74.5 6.5 ;
      RECT 73.5 31.5 74.5 32.5 ;
      RECT 73.5 33.5 74.5 34.5 ;
      RECT 69.5 5.5 70.5 6.5 ;
      RECT 69.5 31.5 70.5 32.5 ;
      RECT 69.5 33.5 70.5 34.5 ;
      RECT 65.5 5.5 66.5 6.5 ;
      RECT 65.5 31.5 66.5 32.5 ;
      RECT 65.5 33.5 66.5 34.5 ;
      RECT 61.5 5.5 62.5 6.5 ;
      RECT 61.5 25.5 62.5 26.5 ;
      RECT 57.5 5.5 58.5 6.5 ;
      RECT 57.5 25.5 58.5 26.5 ;
      RECT 53.5 5.5 54.5 6.5 ;
      RECT 53.5 31.5 54.5 32.5 ;
      RECT 53.5 33.5 54.5 34.5 ;
      RECT 49.5 5.5 50.5 6.5 ;
      RECT 49.5 31.5 50.5 32.5 ;
      RECT 49.5 33.5 50.5 34.5 ;
      RECT 45.5 5.5 46.5 6.5 ;
      RECT 45.5 17.5 46.5 18.5 ;
      RECT 45.5 31.5 46.5 32.5 ;
      RECT 45.5 33.5 46.5 34.5 ;
      RECT 41.5 5.5 42.5 6.5 ;
      RECT 41.5 31.5 42.5 32.5 ;
      RECT 41.5 33.5 42.5 34.5 ;
      RECT 37.5 5.5 38.5 6.5 ;
      RECT 37.5 13.5 38.5 14.5 ;
      RECT 37.5 31.5 38.5 32.5 ;
      RECT 37.5 33.5 38.5 34.5 ;
      RECT 33.5 5.5 34.5 6.5 ;
      RECT 33.5 31.5 34.5 32.5 ;
      RECT 33.5 33.5 34.5 34.5 ;
      RECT 29.5 5.5 30.5 6.5 ;
      RECT 29.5 9.5 30.5 10.5 ;
      RECT 29.5 31.5 30.5 32.5 ;
      RECT 29.5 33.5 30.5 34.5 ;
      RECT 25.5 5.5 26.5 6.5 ;
      RECT 25.5 31.5 26.5 32.5 ;
      RECT 25.5 33.5 26.5 34.5 ;
      RECT 21.5 9.5 22.5 10.5 ;
      RECT 21.5 31.5 22.5 32.5 ;
      RECT 21.5 33.5 22.5 34.5 ;
      RECT 17.5 9.5 18.5 10.5 ;
      RECT 17.5 13.5 18.5 14.5 ;
      RECT 17.5 31.5 18.5 32.5 ;
      RECT 17.5 33.5 18.5 34.5 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 9.5 14.5 10.5 ;
      RECT 13.5 17.5 14.5 18.5 ;
      RECT 13.5 25.5 14.5 26.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 9.5 10.5 10.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 21.5 6.5 22.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END DFFRX1

MACRO DFFSRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRX1 0 0 ;
  SIZE 224 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 224 43 ;
        RECT 217.5 33 221.5 43 ;
        RECT 209.5 33 213.5 43 ;
        RECT 201.5 33 205.5 43 ;
        RECT 178.5 33 182.5 43 ;
        RECT 170.5 33 174.5 43 ;
        RECT 162.5 33 166.5 43 ;
        RECT 149.5 33 153.5 43 ;
        RECT 141.5 33 145.5 43 ;
        RECT 133.5 33 137.5 43 ;
        RECT 110.5 33 114.5 43 ;
        RECT 102.5 33 106.5 43 ;
        RECT 94.5 33 98.5 43 ;
        RECT 81.5 33 85.5 43 ;
        RECT 73.5 33 77.5 43 ;
        RECT 65.5 33 69.5 43 ;
        RECT 42.5 33 46.5 43 ;
        RECT 34.5 33 38.5 43 ;
        RECT 26.5 33 30.5 43 ;
        RECT 17 27 19 43 ;
        RECT 13 27 15 43 ;
        RECT 1 27 3 43 ;
    END
  END VDD!
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 17 13 107 15 ;
        RECT 17 13 19 19 ;
    END
  END SN
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 224 3 ;
        RECT 217 -3 219 7 ;
        RECT 165 -3 167 7 ;
        RECT 149 -3 151 7 ;
        RECT 97 -3 99 7 ;
        RECT 81 -3 83 7 ;
        RECT 29 -3 31 7 ;
        RECT 9 -3 11 7 ;
        RECT 1 -3 3 7 ;
    END
  END VSS!
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9 9 175 11 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 209 21 211 27 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 117 13 123 15 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 125 13 131 15 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 13 3 19 ;
    END
  END RN
  OBS
    LAYER Metal1 ;
      RECT 193 29 221.5 31 ;
      RECT 193 25 195 31 ;
      RECT 37 25 195 27 ;
      RECT 21 21 23 31 ;
      RECT 9 21 11 31 ;
      RECT 9 21 27 23 ;
      RECT 25 17 27 23 ;
      RECT 25 17 219 19 ;
      RECT 5 5 7 31 ;
      RECT 5 17 11 19 ;
      RECT 209 5 215 7 ;
      RECT 201 5 207 7 ;
      RECT 193 5 199 7 ;
      RECT 185 5 191 7 ;
      RECT 157 29 191 31 ;
      RECT 177 5 183 7 ;
      RECT 169 5 175 7 ;
      RECT 97 21 167 23 ;
      RECT 125 29 153.5 31 ;
      RECT 141 5 147 7 ;
      RECT 133 5 139 7 ;
      RECT 125 5 131 7 ;
      RECT 117 5 123 7 ;
      RECT 94.5 29 123 31 ;
      RECT 109 5 115 7 ;
      RECT 101 5 107 7 ;
      RECT 57 29 91 31 ;
      RECT 73 5 79 7 ;
      RECT 65 5 71 7 ;
      RECT 57 5 63 7 ;
      RECT 49 5 55 7 ;
      RECT 26.5 29 55 31 ;
      RECT 41 5 47 7 ;
      RECT 33 5 39 7 ;
      RECT 21 5 27 7 ;
      RECT 13 5 19 7 ;
    LAYER Via1 ;
      RECT 220 29.5 221 30.5 ;
      RECT 220 33.5 221 34.5 ;
      RECT 218 29.5 219 30.5 ;
      RECT 218 33.5 219 34.5 ;
      RECT 217.5 5.5 218.5 6.5 ;
      RECT 217.5 17.5 218.5 18.5 ;
      RECT 213.5 5.5 214.5 6.5 ;
      RECT 212 29.5 213 30.5 ;
      RECT 212 33.5 213 34.5 ;
      RECT 210 29.5 211 30.5 ;
      RECT 210 33.5 211 34.5 ;
      RECT 209.5 5.5 210.5 6.5 ;
      RECT 209.5 25.5 210.5 26.5 ;
      RECT 205.5 5.5 206.5 6.5 ;
      RECT 204 29.5 205 30.5 ;
      RECT 204 33.5 205 34.5 ;
      RECT 202 29.5 203 30.5 ;
      RECT 202 33.5 203 34.5 ;
      RECT 201.5 5.5 202.5 6.5 ;
      RECT 197.5 5.5 198.5 6.5 ;
      RECT 193.5 5.5 194.5 6.5 ;
      RECT 193.5 25.5 194.5 26.5 ;
      RECT 189.5 5.5 190.5 6.5 ;
      RECT 189.5 29.5 190.5 30.5 ;
      RECT 185.5 5.5 186.5 6.5 ;
      RECT 181.5 5.5 182.5 6.5 ;
      RECT 181.5 25.5 182.5 26.5 ;
      RECT 181 29.5 182 30.5 ;
      RECT 181 33.5 182 34.5 ;
      RECT 179 29.5 180 30.5 ;
      RECT 179 33.5 180 34.5 ;
      RECT 177.5 5.5 178.5 6.5 ;
      RECT 173.5 5.5 174.5 6.5 ;
      RECT 173.5 9.5 174.5 10.5 ;
      RECT 173 29.5 174 30.5 ;
      RECT 173 33.5 174 34.5 ;
      RECT 171 29.5 172 30.5 ;
      RECT 171 33.5 172 34.5 ;
      RECT 169.5 5.5 170.5 6.5 ;
      RECT 165.5 5.5 166.5 6.5 ;
      RECT 165.5 21.5 166.5 22.5 ;
      RECT 165 29.5 166 30.5 ;
      RECT 165 33.5 166 34.5 ;
      RECT 163 29.5 164 30.5 ;
      RECT 163 33.5 164 34.5 ;
      RECT 157.5 29.5 158.5 30.5 ;
      RECT 152 29.5 153 30.5 ;
      RECT 152 33.5 153 34.5 ;
      RECT 150 29.5 151 30.5 ;
      RECT 150 33.5 151 34.5 ;
      RECT 149.5 5.5 150.5 6.5 ;
      RECT 145.5 5.5 146.5 6.5 ;
      RECT 144 29.5 145 30.5 ;
      RECT 144 33.5 145 34.5 ;
      RECT 142 29.5 143 30.5 ;
      RECT 142 33.5 143 34.5 ;
      RECT 141.5 5.5 142.5 6.5 ;
      RECT 141.5 17.5 142.5 18.5 ;
      RECT 137.5 5.5 138.5 6.5 ;
      RECT 136 29.5 137 30.5 ;
      RECT 136 33.5 137 34.5 ;
      RECT 134 29.5 135 30.5 ;
      RECT 134 33.5 135 34.5 ;
      RECT 133.5 5.5 134.5 6.5 ;
      RECT 129.5 5.5 130.5 6.5 ;
      RECT 125.5 5.5 126.5 6.5 ;
      RECT 125.5 13.5 126.5 14.5 ;
      RECT 125.5 29.5 126.5 30.5 ;
      RECT 121.5 5.5 122.5 6.5 ;
      RECT 121.5 13.5 122.5 14.5 ;
      RECT 121.5 29.5 122.5 30.5 ;
      RECT 117.5 5.5 118.5 6.5 ;
      RECT 113.5 5.5 114.5 6.5 ;
      RECT 113 29.5 114 30.5 ;
      RECT 113 33.5 114 34.5 ;
      RECT 111 29.5 112 30.5 ;
      RECT 111 33.5 112 34.5 ;
      RECT 109.5 5.5 110.5 6.5 ;
      RECT 105.5 5.5 106.5 6.5 ;
      RECT 105.5 13.5 106.5 14.5 ;
      RECT 105 29.5 106 30.5 ;
      RECT 105 33.5 106 34.5 ;
      RECT 103 29.5 104 30.5 ;
      RECT 103 33.5 104 34.5 ;
      RECT 101.5 5.5 102.5 6.5 ;
      RECT 97.5 5.5 98.5 6.5 ;
      RECT 97.5 21.5 98.5 22.5 ;
      RECT 97 29.5 98 30.5 ;
      RECT 97 33.5 98 34.5 ;
      RECT 95 29.5 96 30.5 ;
      RECT 95 33.5 96 34.5 ;
      RECT 89.5 29.5 90.5 30.5 ;
      RECT 84 29.5 85 30.5 ;
      RECT 84 33.5 85 34.5 ;
      RECT 82 29.5 83 30.5 ;
      RECT 82 33.5 83 34.5 ;
      RECT 81.5 5.5 82.5 6.5 ;
      RECT 81.5 17.5 82.5 18.5 ;
      RECT 77.5 5.5 78.5 6.5 ;
      RECT 76 29.5 77 30.5 ;
      RECT 76 33.5 77 34.5 ;
      RECT 74 29.5 75 30.5 ;
      RECT 74 33.5 75 34.5 ;
      RECT 73.5 5.5 74.5 6.5 ;
      RECT 73.5 9.5 74.5 10.5 ;
      RECT 69.5 5.5 70.5 6.5 ;
      RECT 68 29.5 69 30.5 ;
      RECT 68 33.5 69 34.5 ;
      RECT 66 29.5 67 30.5 ;
      RECT 66 33.5 67 34.5 ;
      RECT 65.5 5.5 66.5 6.5 ;
      RECT 61.5 5.5 62.5 6.5 ;
      RECT 57.5 5.5 58.5 6.5 ;
      RECT 57.5 29.5 58.5 30.5 ;
      RECT 53.5 5.5 54.5 6.5 ;
      RECT 53.5 29.5 54.5 30.5 ;
      RECT 49.5 5.5 50.5 6.5 ;
      RECT 45.5 5.5 46.5 6.5 ;
      RECT 45 29.5 46 30.5 ;
      RECT 45 33.5 46 34.5 ;
      RECT 43 29.5 44 30.5 ;
      RECT 43 33.5 44 34.5 ;
      RECT 41.5 5.5 42.5 6.5 ;
      RECT 37.5 5.5 38.5 6.5 ;
      RECT 37.5 25.5 38.5 26.5 ;
      RECT 37 29.5 38 30.5 ;
      RECT 37 33.5 38 34.5 ;
      RECT 35 29.5 36 30.5 ;
      RECT 35 33.5 36 34.5 ;
      RECT 33.5 5.5 34.5 6.5 ;
      RECT 33.5 13.5 34.5 14.5 ;
      RECT 29.5 5.5 30.5 6.5 ;
      RECT 29 29.5 30 30.5 ;
      RECT 29 33.5 30 34.5 ;
      RECT 27 29.5 28 30.5 ;
      RECT 27 33.5 28 34.5 ;
      RECT 25.5 5.5 26.5 6.5 ;
      RECT 25.5 17.5 26.5 18.5 ;
      RECT 21.5 5.5 22.5 6.5 ;
      RECT 21.5 27.5 22.5 28.5 ;
      RECT 21.5 29.5 22.5 30.5 ;
      RECT 17.5 5.5 18.5 6.5 ;
      RECT 17.5 17.5 18.5 18.5 ;
      RECT 17.5 27.5 18.5 28.5 ;
      RECT 17.5 29.5 18.5 30.5 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 27.5 14.5 28.5 ;
      RECT 13.5 29.5 14.5 30.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 17.5 10.5 18.5 ;
      RECT 9.5 27.5 10.5 28.5 ;
      RECT 9.5 29.5 10.5 30.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 27.5 6.5 28.5 ;
      RECT 5.5 29.5 6.5 30.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 13.5 2.5 14.5 ;
      RECT 1.5 27.5 2.5 28.5 ;
      RECT 1.5 29.5 2.5 30.5 ;
  END
END DFFSRX1

MACRO DFFSX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSX1 0 0 ;
  SIZE 128 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 128 43 ;
        RECT 125 31 127 43 ;
        RECT 113 31 115 43 ;
        RECT 109 31 111 43 ;
        RECT 101 31 103 43 ;
        RECT 93 31 95 43 ;
        RECT 85 31 87 43 ;
        RECT 73 31 75 43 ;
        RECT 61 31 63 43 ;
        RECT 53 31 55 43 ;
        RECT 41 31 43 43 ;
        RECT 33 31 35 43 ;
        RECT 25 31 27 43 ;
        RECT 21 31 23 43 ;
        RECT 13 31 15 43 ;
        RECT 5 31 7 43 ;
    END
  END VDD!
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5 13 51 15 ;
    END
  END SN
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 128 3 ;
        RECT 125 -3 127 11 ;
        RECT 89 -3 91 7 ;
        RECT 85 -3 87 7 ;
        RECT 41 -3 43 7 ;
        RECT 37 -3 39 7 ;
        RECT 1 -3 3 7 ;
    END
  END VSS!
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 37 9 99 11 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 125 13 127 19 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 61 13 67 15 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 69 13 75 15 ;
    END
  END QN
  OBS
    LAYER Metal1 ;
      RECT 117 31 123 35 ;
      RECT 117 17 119 35 ;
      RECT 13 17 119 19 ;
      RECT 113 9 115 19 ;
      RECT 109 5 111 11 ;
      RECT 109 5 115 7 ;
      RECT 105 25 107 35 ;
      RECT 97 25 99 35 ;
      RECT 89 25 91 35 ;
      RECT 85 25 115 27 ;
      RECT 101 9 107 11 ;
      RECT 101 5 103 11 ;
      RECT 77 31 83 35 ;
      RECT 77 25 79 35 ;
      RECT 69 25 79 27 ;
      RECT 57 25 59 35 ;
      RECT 45 31 51 35 ;
      RECT 49 25 51 35 ;
      RECT 49 25 67 27 ;
      RECT 37 25 39 35 ;
      RECT 29 25 31 35 ;
      RECT 21 25 43 27 ;
      RECT 29 9 35 11 ;
      RECT 33 5 35 11 ;
      RECT 25 5 27 11 ;
      RECT 21 5 27 7 ;
      RECT 17 21 19 35 ;
      RECT 9 21 11 35 ;
      RECT 1 21 3 35 ;
      RECT 1 21 27 23 ;
      RECT 117 9 123 11 ;
      RECT 93 5 99 7 ;
      RECT 45 21 91 23 ;
      RECT 77 5 83 7 ;
      RECT 69 5 75 7 ;
      RECT 61 5 67 7 ;
      RECT 53 5 59 7 ;
      RECT 45 5 51 7 ;
      RECT 17 9 23 11 ;
      RECT 13 5 15 11 ;
      RECT 5 5 11 7 ;
    LAYER Via1 ;
      RECT 125.5 9.5 126.5 10.5 ;
      RECT 125.5 17.5 126.5 18.5 ;
      RECT 125.5 31.5 126.5 32.5 ;
      RECT 125.5 33.5 126.5 34.5 ;
      RECT 121.5 9.5 122.5 10.5 ;
      RECT 121.5 31.5 122.5 32.5 ;
      RECT 121.5 33.5 122.5 34.5 ;
      RECT 117.5 9.5 118.5 10.5 ;
      RECT 117.5 31.5 118.5 32.5 ;
      RECT 117.5 33.5 118.5 34.5 ;
      RECT 113.5 5.5 114.5 6.5 ;
      RECT 113.5 9.5 114.5 10.5 ;
      RECT 113.5 25.5 114.5 26.5 ;
      RECT 113.5 31.5 114.5 32.5 ;
      RECT 113.5 33.5 114.5 34.5 ;
      RECT 109.5 9.5 110.5 10.5 ;
      RECT 109.5 31.5 110.5 32.5 ;
      RECT 109.5 33.5 110.5 34.5 ;
      RECT 105.5 9.5 106.5 10.5 ;
      RECT 105.5 17.5 106.5 18.5 ;
      RECT 105.5 31.5 106.5 32.5 ;
      RECT 105.5 33.5 106.5 34.5 ;
      RECT 101.5 5.5 102.5 6.5 ;
      RECT 101.5 31.5 102.5 32.5 ;
      RECT 101.5 33.5 102.5 34.5 ;
      RECT 97.5 5.5 98.5 6.5 ;
      RECT 97.5 9.5 98.5 10.5 ;
      RECT 97.5 31.5 98.5 32.5 ;
      RECT 97.5 33.5 98.5 34.5 ;
      RECT 93.5 5.5 94.5 6.5 ;
      RECT 93.5 31.5 94.5 32.5 ;
      RECT 93.5 33.5 94.5 34.5 ;
      RECT 89.5 5.5 90.5 6.5 ;
      RECT 89.5 21.5 90.5 22.5 ;
      RECT 89.5 31.5 90.5 32.5 ;
      RECT 89.5 33.5 90.5 34.5 ;
      RECT 85.5 5.5 86.5 6.5 ;
      RECT 85.5 25.5 86.5 26.5 ;
      RECT 85.5 31.5 86.5 32.5 ;
      RECT 85.5 33.5 86.5 34.5 ;
      RECT 81.5 5.5 82.5 6.5 ;
      RECT 81.5 31.5 82.5 32.5 ;
      RECT 81.5 33.5 82.5 34.5 ;
      RECT 77.5 5.5 78.5 6.5 ;
      RECT 77.5 31.5 78.5 32.5 ;
      RECT 77.5 33.5 78.5 34.5 ;
      RECT 73.5 5.5 74.5 6.5 ;
      RECT 73.5 31.5 74.5 32.5 ;
      RECT 73.5 33.5 74.5 34.5 ;
      RECT 69.5 5.5 70.5 6.5 ;
      RECT 69.5 13.5 70.5 14.5 ;
      RECT 69.5 25.5 70.5 26.5 ;
      RECT 65.5 5.5 66.5 6.5 ;
      RECT 65.5 13.5 66.5 14.5 ;
      RECT 65.5 25.5 66.5 26.5 ;
      RECT 61.5 5.5 62.5 6.5 ;
      RECT 61.5 31.5 62.5 32.5 ;
      RECT 61.5 33.5 62.5 34.5 ;
      RECT 57.5 5.5 58.5 6.5 ;
      RECT 57.5 31.5 58.5 32.5 ;
      RECT 57.5 33.5 58.5 34.5 ;
      RECT 53.5 5.5 54.5 6.5 ;
      RECT 53.5 31.5 54.5 32.5 ;
      RECT 53.5 33.5 54.5 34.5 ;
      RECT 49.5 5.5 50.5 6.5 ;
      RECT 49.5 13.5 50.5 14.5 ;
      RECT 49.5 31.5 50.5 32.5 ;
      RECT 49.5 33.5 50.5 34.5 ;
      RECT 45.5 5.5 46.5 6.5 ;
      RECT 45.5 21.5 46.5 22.5 ;
      RECT 45.5 31.5 46.5 32.5 ;
      RECT 45.5 33.5 46.5 34.5 ;
      RECT 41.5 5.5 42.5 6.5 ;
      RECT 41.5 25.5 42.5 26.5 ;
      RECT 41.5 31.5 42.5 32.5 ;
      RECT 41.5 33.5 42.5 34.5 ;
      RECT 37.5 5.5 38.5 6.5 ;
      RECT 37.5 9.5 38.5 10.5 ;
      RECT 37.5 31.5 38.5 32.5 ;
      RECT 37.5 33.5 38.5 34.5 ;
      RECT 33.5 5.5 34.5 6.5 ;
      RECT 33.5 31.5 34.5 32.5 ;
      RECT 33.5 33.5 34.5 34.5 ;
      RECT 29.5 9.5 30.5 10.5 ;
      RECT 29.5 31.5 30.5 32.5 ;
      RECT 29.5 33.5 30.5 34.5 ;
      RECT 25.5 9.5 26.5 10.5 ;
      RECT 25.5 21.5 26.5 22.5 ;
      RECT 25.5 31.5 26.5 32.5 ;
      RECT 25.5 33.5 26.5 34.5 ;
      RECT 21.5 5.5 22.5 6.5 ;
      RECT 21.5 9.5 22.5 10.5 ;
      RECT 21.5 25.5 22.5 26.5 ;
      RECT 21.5 31.5 22.5 32.5 ;
      RECT 21.5 33.5 22.5 34.5 ;
      RECT 17.5 9.5 18.5 10.5 ;
      RECT 17.5 31.5 18.5 32.5 ;
      RECT 17.5 33.5 18.5 34.5 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 9.5 14.5 10.5 ;
      RECT 13.5 17.5 14.5 18.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 13.5 6.5 14.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END DFFSX1

MACRO DFFX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFX1 0 0 ;
  SIZE 108 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 108 43 ;
        RECT 101 27 103 43 ;
        RECT 97 27 99 43 ;
        RECT 85 31 87 43 ;
        RECT 81 31 83 43 ;
        RECT 69 31 71 43 ;
        RECT 65 31 67 43 ;
        RECT 57 31 59 43 ;
        RECT 41 31 43 43 ;
        RECT 33 31 35 43 ;
        RECT 29 31 31 43 ;
        RECT 17 31 19 43 ;
        RECT 13 31 15 43 ;
        RECT 1 31 3 43 ;
    END
  END VDD!
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 108 3 ;
        RECT 105 -3 107 11 ;
        RECT 69 -3 71 7 ;
        RECT 65 -3 67 7 ;
        RECT 33 -3 35 7 ;
        RECT 29 -3 31 7 ;
        RECT 1 -3 3 7 ;
    END
  END VSS!
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 29 13 79 15 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 105 13 107 19 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 45 31 51 35 ;
        RECT 45 25 47 35 ;
        RECT 37 25 47 27 ;
        RECT 37 25 39 35 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 61 25 63 35 ;
        RECT 49 25 63 27 ;
        RECT 53 25 55 35 ;
    END
  END QN
  OBS
    LAYER Metal1 ;
      RECT 105 21 107 31 ;
      RECT 93 9 95 31 ;
      RECT 93 21 107 23 ;
      RECT 5 17 95 19 ;
      RECT 89 33 95 35 ;
      RECT 73 31 79 35 ;
      RECT 89 25 91 35 ;
      RECT 73 25 75 35 ;
      RECT 65 25 91 27 ;
      RECT 21 31 27 35 ;
      RECT 25 21 27 35 ;
      RECT 13 21 75 23 ;
      RECT 57 5 59 11 ;
      RECT 57 5 63 7 ;
      RECT 21 5 23 11 ;
      RECT 21 5 27 7 ;
      RECT 5 31 11 35 ;
      RECT 9 25 11 35 ;
      RECT 9 25 19 27 ;
      RECT 97 9 103 11 ;
      RECT 89 5 95 7 ;
      RECT 81 5 87 7 ;
      RECT 73 5 79 7 ;
      RECT 45 5 55 7 ;
      RECT 45 9 55 11 ;
      RECT 37 5 43 7 ;
      RECT 13 5 19 7 ;
      RECT 13 9 19 11 ;
      RECT 5 5 11 7 ;
    LAYER Via1 ;
      RECT 105.5 9.5 106.5 10.5 ;
      RECT 105.5 13.5 106.5 14.5 ;
      RECT 105.5 27.5 106.5 28.5 ;
      RECT 105.5 29.5 106.5 30.5 ;
      RECT 101.5 9.5 102.5 10.5 ;
      RECT 101.5 27.5 102.5 28.5 ;
      RECT 101.5 29.5 102.5 30.5 ;
      RECT 97.5 9.5 98.5 10.5 ;
      RECT 97.5 27.5 98.5 28.5 ;
      RECT 97.5 29.5 98.5 30.5 ;
      RECT 93.5 5.5 94.5 6.5 ;
      RECT 93.5 9.5 94.5 10.5 ;
      RECT 93.5 27.5 94.5 28.5 ;
      RECT 93.5 29.5 94.5 30.5 ;
      RECT 93.5 33.5 94.5 34.5 ;
      RECT 89.5 5.5 90.5 6.5 ;
      RECT 89.5 31.5 90.5 32.5 ;
      RECT 89.5 33.5 90.5 34.5 ;
      RECT 85.5 5.5 86.5 6.5 ;
      RECT 85.5 17.5 86.5 18.5 ;
      RECT 85.5 31.5 86.5 32.5 ;
      RECT 85.5 33.5 86.5 34.5 ;
      RECT 81.5 5.5 82.5 6.5 ;
      RECT 81.5 31.5 82.5 32.5 ;
      RECT 81.5 33.5 82.5 34.5 ;
      RECT 77.5 5.5 78.5 6.5 ;
      RECT 77.5 13.5 78.5 14.5 ;
      RECT 77.5 31.5 78.5 32.5 ;
      RECT 77.5 33.5 78.5 34.5 ;
      RECT 73.5 5.5 74.5 6.5 ;
      RECT 73.5 31.5 74.5 32.5 ;
      RECT 73.5 33.5 74.5 34.5 ;
      RECT 69.5 5.5 70.5 6.5 ;
      RECT 69.5 21.5 70.5 22.5 ;
      RECT 69.5 31.5 70.5 32.5 ;
      RECT 69.5 33.5 70.5 34.5 ;
      RECT 65.5 5.5 66.5 6.5 ;
      RECT 65.5 25.5 66.5 26.5 ;
      RECT 65.5 31.5 66.5 32.5 ;
      RECT 65.5 33.5 66.5 34.5 ;
      RECT 61.5 5.5 62.5 6.5 ;
      RECT 61.5 31.5 62.5 32.5 ;
      RECT 61.5 33.5 62.5 34.5 ;
      RECT 57.5 9.5 58.5 10.5 ;
      RECT 57.5 31.5 58.5 32.5 ;
      RECT 57.5 33.5 58.5 34.5 ;
      RECT 53.5 5.5 54.5 6.5 ;
      RECT 53.5 9.5 54.5 10.5 ;
      RECT 53.5 31.5 54.5 32.5 ;
      RECT 53.5 33.5 54.5 34.5 ;
      RECT 49.5 25.5 50.5 26.5 ;
      RECT 49.5 31.5 50.5 32.5 ;
      RECT 49.5 33.5 50.5 34.5 ;
      RECT 45.5 5.5 46.5 6.5 ;
      RECT 45.5 9.5 46.5 10.5 ;
      RECT 45.5 31.5 46.5 32.5 ;
      RECT 45.5 33.5 46.5 34.5 ;
      RECT 41.5 5.5 42.5 6.5 ;
      RECT 41.5 31.5 42.5 32.5 ;
      RECT 41.5 33.5 42.5 34.5 ;
      RECT 37.5 5.5 38.5 6.5 ;
      RECT 37.5 31.5 38.5 32.5 ;
      RECT 37.5 33.5 38.5 34.5 ;
      RECT 33.5 5.5 34.5 6.5 ;
      RECT 33.5 21.5 34.5 22.5 ;
      RECT 33.5 31.5 34.5 32.5 ;
      RECT 33.5 33.5 34.5 34.5 ;
      RECT 29.5 5.5 30.5 6.5 ;
      RECT 29.5 13.5 30.5 14.5 ;
      RECT 29.5 31.5 30.5 32.5 ;
      RECT 29.5 33.5 30.5 34.5 ;
      RECT 25.5 5.5 26.5 6.5 ;
      RECT 25.5 31.5 26.5 32.5 ;
      RECT 25.5 33.5 26.5 34.5 ;
      RECT 21.5 9.5 22.5 10.5 ;
      RECT 21.5 31.5 22.5 32.5 ;
      RECT 21.5 33.5 22.5 34.5 ;
      RECT 17.5 5.5 18.5 6.5 ;
      RECT 17.5 9.5 18.5 10.5 ;
      RECT 17.5 25.5 18.5 26.5 ;
      RECT 17.5 31.5 18.5 32.5 ;
      RECT 17.5 33.5 18.5 34.5 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 9.5 14.5 10.5 ;
      RECT 13.5 21.5 14.5 22.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 17.5 6.5 18.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END DFFX1

MACRO FILL1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL1 0 0 ;
  SIZE 4 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 4 43 ;
    END
  END VDD!
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 4 3 ;
    END
  END VSS!
END FILL1

MACRO FILL2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL2 0 0 ;
  SIZE 8 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 8 43 ;
    END
  END VDD!
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 8 3 ;
    END
  END VSS!
END FILL2

MACRO FILL3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL3 0 0 ;
  SIZE 16 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 16 43 ;
    END
  END VDD!
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 16 3 ;
    END
  END VSS!
END FILL3

MACRO FILL4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL4 0 0 ;
  SIZE 32 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 32 43 ;
    END
  END VDD!
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 32 3 ;
    END
  END VSS!
END FILL4

MACRO INVX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX1 0 0 ;
  SIZE 8 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5 5 7 35 ;
    END
  END Y
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 8 43 ;
        RECT 1 31 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 17 3 23 ;
    END
  END A
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 8 3 ;
        RECT 1 -3 3 7 ;
    END
  END VSS!
  OBS
    LAYER Via1 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 21.5 2.5 22.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END INVX1

MACRO INVX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX2 0 0 ;
  SIZE 8 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5 5 7 35 ;
    END
  END Y
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 8 43 ;
        RECT 1 27 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 13 3 19 ;
    END
  END A
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 8 3 ;
        RECT 1 -3 3 9 ;
    END
  END VSS!
  OBS
    LAYER Via1 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 7.5 6.5 8.5 ;
      RECT 5.5 27.5 6.5 28.5 ;
      RECT 5.5 29.5 6.5 30.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 7.5 2.5 8.5 ;
      RECT 1.5 17.5 2.5 18.5 ;
      RECT 1.5 27.5 2.5 28.5 ;
      RECT 1.5 29.5 2.5 30.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END INVX2

MACRO INVX3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX3 0 0 ;
  SIZE 8 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5 5 7 35 ;
    END
  END Y
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 8 43 ;
        RECT 1 23 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 13 3 19 ;
    END
  END A
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 8 3 ;
        RECT 1 -3 3 11 ;
    END
  END VSS!
  OBS
    LAYER Via1 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 7.5 6.5 8.5 ;
      RECT 5.5 9.5 6.5 10.5 ;
      RECT 5.5 23.5 6.5 24.5 ;
      RECT 5.5 25.5 6.5 26.5 ;
      RECT 5.5 27.5 6.5 28.5 ;
      RECT 5.5 29.5 6.5 30.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 7.5 2.5 8.5 ;
      RECT 1.5 9.5 2.5 10.5 ;
      RECT 1.5 13.5 2.5 14.5 ;
      RECT 1.5 23.5 2.5 24.5 ;
      RECT 1.5 25.5 2.5 26.5 ;
      RECT 1.5 27.5 2.5 28.5 ;
      RECT 1.5 29.5 2.5 30.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END INVX3

MACRO INVX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX4 0 0 ;
  SIZE 12 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5 5 7 35 ;
    END
  END Y
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 12 43 ;
        RECT 9 27 11 43 ;
        RECT 1 27 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 13 3 19 ;
    END
  END A
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 12 3 ;
        RECT 9 -3 11 9 ;
        RECT 1 -3 3 9 ;
    END
  END VSS!
  OBS
    LAYER Via1 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 7.5 10.5 8.5 ;
      RECT 9.5 27.5 10.5 28.5 ;
      RECT 9.5 29.5 10.5 30.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 7.5 6.5 8.5 ;
      RECT 5.5 27.5 6.5 28.5 ;
      RECT 5.5 29.5 6.5 30.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 7.5 2.5 8.5 ;
      RECT 1.5 17.5 2.5 18.5 ;
      RECT 1.5 27.5 2.5 28.5 ;
      RECT 1.5 29.5 2.5 30.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END INVX4

MACRO MX2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX2X1 0 0 ;
  SIZE 48 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 48 43 ;
        RECT 41 27 43 43 ;
        RECT 37 27 39 43 ;
        RECT 9 27 11 43 ;
        RECT 1 27 3 43 ;
    END
  END VDD!
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 13 3 19 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 45 9 47 31 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 48 3 ;
        RECT 41 -3 43 11 ;
        RECT 37 -3 39 11 ;
        RECT 9 -3 11 11 ;
        RECT 1 -3 3 11 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 33 13 35 19 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 13 21 19 23 ;
    END
  END B
  OBS
    LAYER Metal1 ;
      RECT 21 27 27 31 ;
      RECT 25 9 27 31 ;
      RECT 25 21 43 23 ;
      RECT 21 9 27 11 ;
      RECT 5 9 7 31 ;
      RECT 5 17 19 19 ;
      RECT 29 9 35 11 ;
      RECT 29 27 35 31 ;
      RECT 13 9 19 11 ;
      RECT 13 27 19 31 ;
    LAYER Via1 ;
      RECT 45.5 9.5 46.5 10.5 ;
      RECT 45.5 27.5 46.5 28.5 ;
      RECT 45.5 29.5 46.5 30.5 ;
      RECT 41.5 9.5 42.5 10.5 ;
      RECT 41.5 21.5 42.5 22.5 ;
      RECT 41.5 27.5 42.5 28.5 ;
      RECT 41.5 29.5 42.5 30.5 ;
      RECT 37.5 9.5 38.5 10.5 ;
      RECT 37.5 27.5 38.5 28.5 ;
      RECT 37.5 29.5 38.5 30.5 ;
      RECT 33.5 9.5 34.5 10.5 ;
      RECT 33.5 13.5 34.5 14.5 ;
      RECT 33.5 27.5 34.5 28.5 ;
      RECT 33.5 29.5 34.5 30.5 ;
      RECT 29.5 9.5 30.5 10.5 ;
      RECT 29.5 27.5 30.5 28.5 ;
      RECT 29.5 29.5 30.5 30.5 ;
      RECT 25.5 9.5 26.5 10.5 ;
      RECT 25.5 27.5 26.5 28.5 ;
      RECT 25.5 29.5 26.5 30.5 ;
      RECT 21.5 9.5 22.5 10.5 ;
      RECT 21.5 27.5 22.5 28.5 ;
      RECT 21.5 29.5 22.5 30.5 ;
      RECT 17.5 9.5 18.5 10.5 ;
      RECT 17.5 17.5 18.5 18.5 ;
      RECT 17.5 27.5 18.5 28.5 ;
      RECT 17.5 29.5 18.5 30.5 ;
      RECT 13.5 9.5 14.5 10.5 ;
      RECT 13.5 21.5 14.5 22.5 ;
      RECT 13.5 27.5 14.5 28.5 ;
      RECT 13.5 29.5 14.5 30.5 ;
      RECT 9.5 9.5 10.5 10.5 ;
      RECT 9.5 27.5 10.5 28.5 ;
      RECT 9.5 29.5 10.5 30.5 ;
      RECT 5.5 9.5 6.5 10.5 ;
      RECT 5.5 27.5 6.5 28.5 ;
      RECT 5.5 29.5 6.5 30.5 ;
      RECT 1.5 9.5 2.5 10.5 ;
      RECT 1.5 17.5 2.5 18.5 ;
      RECT 1.5 27.5 2.5 28.5 ;
      RECT 1.5 29.5 2.5 30.5 ;
  END
END MX2X1

MACRO MX4X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX4X1 0 0 ;
  SIZE 140 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 140 43 ;
        RECT 133 31 135 43 ;
        RECT 105 33 109 43 ;
        RECT 69 29 71 43 ;
        RECT 37 33 41 43 ;
        RECT 1 31 3 43 ;
    END
  END VDD!
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 21 127 23 ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 41 13 111 15 ;
    END
  END S1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 137 5 139 35 ;
    END
  END Y
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 113 5 119 7 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 101 5 107 7 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 45 5 51 7 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 33 5 39 7 ;
    END
  END A
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 140 3 ;
        RECT 133 -3 135 7 ;
        RECT 109 -3 111 7 ;
        RECT 69 -3 71 11 ;
        RECT 41 -3 43 7 ;
        RECT 1 -3 3 7 ;
    END
  END VSS!
  OBS
    LAYER Metal1 ;
      RECT 127 29 131 31 ;
      RECT 129 9 131 31 ;
      RECT 13 17 135 19 ;
      RECT 121 5 131 7 ;
      RECT 113 33 131 35 ;
      RECT 9 25 127 27 ;
      RECT 97 9 123 11 ;
      RECT 95 29 117 31 ;
      RECT 89 5 99 7 ;
      RECT 85 33 99 35 ;
      RECT 81 9 91 11 ;
      RECT 81 29 89 31 ;
      RECT 73 9 79 11 ;
      RECT 73 29 79 33 ;
      RECT 61 9 67 11 ;
      RECT 57 29 67 31 ;
      RECT 53 5 63 7 ;
      RECT 45 33 61 35 ;
      RECT 29 9 55 11 ;
      RECT 27 29 49 31 ;
      RECT 21 5 31 7 ;
      RECT 17 33 31 35 ;
      RECT 13 9 23 11 ;
      RECT 13 29 21 31 ;
      RECT 5 5 11 7 ;
      RECT 5 31 11 35 ;
    LAYER Via1 ;
      RECT 137.5 5.5 138.5 6.5 ;
      RECT 137.5 31.5 138.5 32.5 ;
      RECT 137.5 33.5 138.5 34.5 ;
      RECT 133.5 5.5 134.5 6.5 ;
      RECT 133.5 17.5 134.5 18.5 ;
      RECT 133.5 31.5 134.5 32.5 ;
      RECT 133.5 33.5 134.5 34.5 ;
      RECT 129.5 5.5 130.5 6.5 ;
      RECT 129.5 9.5 130.5 10.5 ;
      RECT 129.5 29.5 130.5 30.5 ;
      RECT 129.5 33.5 130.5 34.5 ;
      RECT 127.5 29.5 128.5 30.5 ;
      RECT 127.5 33.5 128.5 34.5 ;
      RECT 125.5 21.5 126.5 22.5 ;
      RECT 125.5 25.5 126.5 26.5 ;
      RECT 121.5 5.5 122.5 6.5 ;
      RECT 121.5 9.5 122.5 10.5 ;
      RECT 117.5 5.5 118.5 6.5 ;
      RECT 115.5 29.5 116.5 30.5 ;
      RECT 115.5 33.5 116.5 34.5 ;
      RECT 113.5 29.5 114.5 30.5 ;
      RECT 113.5 33.5 114.5 34.5 ;
      RECT 109.5 5.5 110.5 6.5 ;
      RECT 109.5 9.5 110.5 10.5 ;
      RECT 109.5 13.5 110.5 14.5 ;
      RECT 107.5 29.5 108.5 30.5 ;
      RECT 107.5 33.5 108.5 34.5 ;
      RECT 105.5 29.5 106.5 30.5 ;
      RECT 105.5 33.5 106.5 34.5 ;
      RECT 101.5 5.5 102.5 6.5 ;
      RECT 97.5 5.5 98.5 6.5 ;
      RECT 97.5 9.5 98.5 10.5 ;
      RECT 97.5 29.5 98.5 30.5 ;
      RECT 97.5 33.5 98.5 34.5 ;
      RECT 95.5 29.5 96.5 30.5 ;
      RECT 95.5 33.5 96.5 34.5 ;
      RECT 89.5 5.5 90.5 6.5 ;
      RECT 89.5 9.5 90.5 10.5 ;
      RECT 89.5 21.5 90.5 22.5 ;
      RECT 87.5 29.5 88.5 30.5 ;
      RECT 87.5 33.5 88.5 34.5 ;
      RECT 85.5 25.5 86.5 26.5 ;
      RECT 85.5 29.5 86.5 30.5 ;
      RECT 85.5 33.5 86.5 34.5 ;
      RECT 81.5 9.5 82.5 10.5 ;
      RECT 81.5 17.5 82.5 18.5 ;
      RECT 81.5 29.5 82.5 30.5 ;
      RECT 77.5 9.5 78.5 10.5 ;
      RECT 77.5 29.5 78.5 30.5 ;
      RECT 77.5 31.5 78.5 32.5 ;
      RECT 73.5 9.5 74.5 10.5 ;
      RECT 73.5 29.5 74.5 30.5 ;
      RECT 73.5 31.5 74.5 32.5 ;
      RECT 69.5 9.5 70.5 10.5 ;
      RECT 69.5 13.5 70.5 14.5 ;
      RECT 69.5 29.5 70.5 30.5 ;
      RECT 69.5 31.5 70.5 32.5 ;
      RECT 65.5 9.5 66.5 10.5 ;
      RECT 65.5 17.5 66.5 18.5 ;
      RECT 65.5 29.5 66.5 30.5 ;
      RECT 61.5 5.5 62.5 6.5 ;
      RECT 61.5 9.5 62.5 10.5 ;
      RECT 59.5 29.5 60.5 30.5 ;
      RECT 59.5 33.5 60.5 34.5 ;
      RECT 57.5 21.5 58.5 22.5 ;
      RECT 57.5 25.5 58.5 26.5 ;
      RECT 57.5 29.5 58.5 30.5 ;
      RECT 57.5 33.5 58.5 34.5 ;
      RECT 53.5 5.5 54.5 6.5 ;
      RECT 53.5 9.5 54.5 10.5 ;
      RECT 49.5 5.5 50.5 6.5 ;
      RECT 47.5 29.5 48.5 30.5 ;
      RECT 47.5 33.5 48.5 34.5 ;
      RECT 45.5 29.5 46.5 30.5 ;
      RECT 45.5 33.5 46.5 34.5 ;
      RECT 41.5 5.5 42.5 6.5 ;
      RECT 41.5 9.5 42.5 10.5 ;
      RECT 41.5 13.5 42.5 14.5 ;
      RECT 39.5 29.5 40.5 30.5 ;
      RECT 39.5 33.5 40.5 34.5 ;
      RECT 37.5 29.5 38.5 30.5 ;
      RECT 37.5 33.5 38.5 34.5 ;
      RECT 33.5 5.5 34.5 6.5 ;
      RECT 29.5 5.5 30.5 6.5 ;
      RECT 29.5 9.5 30.5 10.5 ;
      RECT 29.5 29.5 30.5 30.5 ;
      RECT 29.5 33.5 30.5 34.5 ;
      RECT 27.5 29.5 28.5 30.5 ;
      RECT 27.5 33.5 28.5 34.5 ;
      RECT 21.5 5.5 22.5 6.5 ;
      RECT 21.5 9.5 22.5 10.5 ;
      RECT 21.5 21.5 22.5 22.5 ;
      RECT 19.5 29.5 20.5 30.5 ;
      RECT 19.5 33.5 20.5 34.5 ;
      RECT 17.5 25.5 18.5 26.5 ;
      RECT 17.5 29.5 18.5 30.5 ;
      RECT 17.5 33.5 18.5 34.5 ;
      RECT 13.5 9.5 14.5 10.5 ;
      RECT 13.5 17.5 14.5 18.5 ;
      RECT 13.5 29.5 14.5 30.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 25.5 10.5 26.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 21.5 2.5 22.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END MX4X1

MACRO NAND2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X1 0 0 ;
  SIZE 16 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9 25 15 27 ;
        RECT 13 5 15 27 ;
        RECT 5 31 11 35 ;
        RECT 9 25 11 35 ;
    END
  END Y
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 16 43 ;
        RECT 13 31 15 43 ;
        RECT 1 31 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 9 3 15 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9 13 11 19 ;
    END
  END B
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 16 3 ;
        RECT 1 -3 3 7 ;
    END
  END VSS!
  OBS
    LAYER Metal1 ;
      RECT 5 5 11 7 ;
    LAYER Via1 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 13.5 10.5 14.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 9.5 2.5 10.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END NAND2X1

MACRO NAND2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X2 0 0 ;
  SIZE 16 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9 21 15 23 ;
        RECT 13 5 15 23 ;
        RECT 5 27 11 35 ;
        RECT 9 21 11 35 ;
    END
  END Y
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 16 43 ;
        RECT 13 27 15 43 ;
        RECT 1 27 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 17 3 23 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5 13 11 15 ;
    END
  END B
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 16 3 ;
        RECT 1 -3 3 9 ;
    END
  END VSS!
  OBS
    LAYER Metal1 ;
      RECT 5 5 11 9 ;
    LAYER Via1 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 7.5 14.5 8.5 ;
      RECT 13.5 27.5 14.5 28.5 ;
      RECT 13.5 29.5 14.5 30.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 7.5 10.5 8.5 ;
      RECT 9.5 13.5 10.5 14.5 ;
      RECT 9.5 27.5 10.5 28.5 ;
      RECT 9.5 29.5 10.5 30.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 7.5 6.5 8.5 ;
      RECT 5.5 27.5 6.5 28.5 ;
      RECT 5.5 29.5 6.5 30.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 7.5 2.5 8.5 ;
      RECT 1.5 17.5 2.5 18.5 ;
      RECT 1.5 27.5 2.5 28.5 ;
      RECT 1.5 29.5 2.5 30.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END NAND2X2

MACRO NAND2X3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X3 0 0 ;
  SIZE 24 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 17 5 19 35 ;
        RECT 5 25 19 27 ;
        RECT 5 25 7 35 ;
    END
  END Y
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 24 43 ;
        RECT 21 29 23 43 ;
        RECT 13 29 15 43 ;
        RECT 9 29 11 43 ;
        RECT 1 29 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 13 7 15 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9 17 15 19 ;
    END
  END B
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 24 3 ;
        RECT 5 -3 7 11 ;
    END
  END VSS!
  OBS
    LAYER Metal1 ;
      RECT 9 5 15 11 ;
    LAYER Via1 ;
      RECT 21.5 29.5 22.5 30.5 ;
      RECT 21.5 31.5 22.5 32.5 ;
      RECT 21.5 33.5 22.5 34.5 ;
      RECT 17.5 5.5 18.5 6.5 ;
      RECT 17.5 7.5 18.5 8.5 ;
      RECT 17.5 9.5 18.5 10.5 ;
      RECT 17.5 29.5 18.5 30.5 ;
      RECT 17.5 31.5 18.5 32.5 ;
      RECT 17.5 33.5 18.5 34.5 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 7.5 14.5 8.5 ;
      RECT 13.5 9.5 14.5 10.5 ;
      RECT 13.5 17.5 14.5 18.5 ;
      RECT 13.5 29.5 14.5 30.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 7.5 10.5 8.5 ;
      RECT 9.5 9.5 10.5 10.5 ;
      RECT 9.5 29.5 10.5 30.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 7.5 6.5 8.5 ;
      RECT 5.5 9.5 6.5 10.5 ;
      RECT 5.5 13.5 6.5 14.5 ;
      RECT 5.5 29.5 6.5 30.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 29.5 2.5 30.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END NAND2X3

MACRO NAND3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X1 0 0 ;
  SIZE 24 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 24 43 ;
        RECT 17 31 19 43 ;
        RECT 9 31 11 43 ;
        RECT 1 31 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 21 3 27 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9 13 11 19 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 17 9 19 15 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 21 5 23 35 ;
        RECT 5 25 23 27 ;
        RECT 13 25 15 35 ;
        RECT 5 25 7 35 ;
    END
  END Y
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 24 3 ;
        RECT 1 -3 3 7 ;
    END
  END VSS!
  OBS
    LAYER Metal1 ;
      RECT 13 5 19 7 ;
      RECT 5 5 11 7 ;
    LAYER Via1 ;
      RECT 21.5 5.5 22.5 6.5 ;
      RECT 21.5 31.5 22.5 32.5 ;
      RECT 21.5 33.5 22.5 34.5 ;
      RECT 17.5 5.5 18.5 6.5 ;
      RECT 17.5 13.5 18.5 14.5 ;
      RECT 17.5 31.5 18.5 32.5 ;
      RECT 17.5 33.5 18.5 34.5 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 13.5 10.5 14.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 21.5 2.5 22.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END NAND3X1

MACRO NAND4X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X1 0 0 ;
  SIZE 32 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 32 43 ;
        RECT 25 31 27 43 ;
        RECT 17 31 19 43 ;
        RECT 9 31 11 43 ;
        RECT 1 31 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 21 3 27 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9 17 15 19 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 17 13 19 19 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 25 9 27 15 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 29 5 31 35 ;
        RECT 5 25 31 27 ;
        RECT 21 25 23 35 ;
        RECT 13 25 15 35 ;
        RECT 5 25 7 35 ;
    END
  END Y
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 32 3 ;
        RECT 1 -3 3 7 ;
    END
  END VSS!
  OBS
    LAYER Metal1 ;
      RECT 21 5 27 7 ;
      RECT 13 5 19 7 ;
      RECT 5 5 11 7 ;
    LAYER Via1 ;
      RECT 29.5 5.5 30.5 6.5 ;
      RECT 29.5 31.5 30.5 32.5 ;
      RECT 29.5 33.5 30.5 34.5 ;
      RECT 25.5 5.5 26.5 6.5 ;
      RECT 25.5 13.5 26.5 14.5 ;
      RECT 25.5 31.5 26.5 32.5 ;
      RECT 25.5 33.5 26.5 34.5 ;
      RECT 21.5 5.5 22.5 6.5 ;
      RECT 21.5 31.5 22.5 32.5 ;
      RECT 21.5 33.5 22.5 34.5 ;
      RECT 17.5 5.5 18.5 6.5 ;
      RECT 17.5 17.5 18.5 18.5 ;
      RECT 17.5 31.5 18.5 32.5 ;
      RECT 17.5 33.5 18.5 34.5 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 17.5 14.5 18.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 25.5 2.5 26.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END NAND4X1

MACRO NOR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X1 0 0 ;
  SIZE 16 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 16 43 ;
        RECT 1 31 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 9 3 15 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5 17 11 19 ;
    END
  END B
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 16 3 ;
        RECT 9 -3 11 7 ;
        RECT 1 -3 3 7 ;
    END
  END VSS!
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 13 5 15 35 ;
        RECT 5 9 15 11 ;
        RECT 5 5 7 11 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 5 31 11 35 ;
    LAYER Via1 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 17.5 10.5 18.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 13.5 2.5 14.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END NOR2X1

MACRO NOR2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X2 0 0 ;
  SIZE 16 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 16 43 ;
        RECT 1 27 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 13 3 19 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5 21 11 23 ;
    END
  END B
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 16 3 ;
        RECT 9 -3 11 9 ;
        RECT 1 -3 3 9 ;
    END
  END VSS!
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 13 5 15 35 ;
        RECT 5 13 15 15 ;
        RECT 5 5 7 15 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 5 27 11 35 ;
    LAYER Via1 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 7.5 14.5 8.5 ;
      RECT 13.5 27.5 14.5 28.5 ;
      RECT 13.5 29.5 14.5 30.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 7.5 10.5 8.5 ;
      RECT 9.5 21.5 10.5 22.5 ;
      RECT 9.5 27.5 10.5 28.5 ;
      RECT 9.5 29.5 10.5 30.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 7.5 6.5 8.5 ;
      RECT 5.5 27.5 6.5 28.5 ;
      RECT 5.5 29.5 6.5 30.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 7.5 2.5 8.5 ;
      RECT 1.5 17.5 2.5 18.5 ;
      RECT 1.5 27.5 2.5 28.5 ;
      RECT 1.5 29.5 2.5 30.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END NOR2X2

MACRO NOR2X3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X3 0 0 ;
  SIZE 24 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 24 43 ;
        RECT 9 29 11 43 ;
        RECT 1 29 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 17 7 19 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9 21 15 23 ;
    END
  END B
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 24 3 ;
        RECT 13 -3 15 11 ;
        RECT 9 -3 11 11 ;
    END
  END VSS!
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 17 5 19 31 ;
        RECT 5 13 19 15 ;
        RECT 5 5 7 15 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 13 33 23 35 ;
      RECT 21 25 23 35 ;
      RECT 5 25 7 35 ;
      RECT 13 25 15 35 ;
      RECT 5 25 15 27 ;
    LAYER Via1 ;
      RECT 21.55 25.5 22.55 26.5 ;
      RECT 21.55 27.5 22.55 28.5 ;
      RECT 21.55 29.5 22.55 30.5 ;
      RECT 17.5 5.5 18.5 6.5 ;
      RECT 17.5 7.5 18.5 8.5 ;
      RECT 17.5 9.5 18.5 10.5 ;
      RECT 17.5 25.5 18.5 26.5 ;
      RECT 17.5 27.5 18.5 28.5 ;
      RECT 17.5 29.5 18.5 30.5 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 7.5 14.5 8.5 ;
      RECT 13.5 9.5 14.5 10.5 ;
      RECT 13.5 21.5 14.5 22.5 ;
      RECT 13.5 25.5 14.5 26.5 ;
      RECT 13.5 27.5 14.5 28.5 ;
      RECT 13.5 29.5 14.5 30.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 7.5 10.5 8.5 ;
      RECT 9.5 9.5 10.5 10.5 ;
      RECT 9.5 29.5 10.5 30.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 7.5 6.5 8.5 ;
      RECT 5.5 9.5 6.5 10.5 ;
      RECT 5.5 17.5 6.5 18.5 ;
      RECT 5.5 29.5 6.5 30.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 29.5 2.5 30.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END NOR2X3

MACRO NOR3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X1 0 0 ;
  SIZE 24 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 24 43 ;
        RECT 1 31 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 9 3 15 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9 17 11 23 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 17 21 19 27 ;
    END
  END C
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 24 3 ;
        RECT 17 -3 19 7 ;
        RECT 9 -3 11 7 ;
        RECT 1 -3 3 7 ;
    END
  END VSS!
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 21 5 23 35 ;
        RECT 5 9 23 11 ;
        RECT 13 5 15 11 ;
        RECT 5 5 7 11 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 13 31 19 35 ;
      RECT 5 31 11 35 ;
    LAYER Via1 ;
      RECT 21.5 5.5 22.5 6.5 ;
      RECT 21.5 31.5 22.5 32.5 ;
      RECT 21.5 33.5 22.5 34.5 ;
      RECT 17.5 5.5 18.5 6.5 ;
      RECT 17.5 21.5 18.5 22.5 ;
      RECT 17.5 31.5 18.5 32.5 ;
      RECT 17.5 33.5 18.5 34.5 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 21.5 10.5 22.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 13.5 2.5 14.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END NOR3X1

MACRO NOR4X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X1 0 0 ;
  SIZE 32 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 32 43 ;
        RECT 1 31 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 9 3 15 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9 17 15 19 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 17 17 19 23 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 25 21 27 27 ;
    END
  END D
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 32 3 ;
        RECT 25 -3 27 7 ;
        RECT 17 -3 19 7 ;
        RECT 9 -3 11 7 ;
        RECT 1 -3 3 7 ;
    END
  END VSS!
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 29 5 31 35 ;
        RECT 5 9 31 11 ;
        RECT 21 5 23 11 ;
        RECT 13 5 15 11 ;
        RECT 5 5 7 11 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 21 31 27 35 ;
      RECT 13 31 19 35 ;
      RECT 5 31 11 35 ;
    LAYER Via1 ;
      RECT 29.5 5.5 30.5 6.5 ;
      RECT 29.5 31.5 30.5 32.5 ;
      RECT 29.5 33.5 30.5 34.5 ;
      RECT 25.5 5.5 26.5 6.5 ;
      RECT 25.5 21.5 26.5 22.5 ;
      RECT 25.5 31.5 26.5 32.5 ;
      RECT 25.5 33.5 26.5 34.5 ;
      RECT 21.5 5.5 22.5 6.5 ;
      RECT 21.5 31.5 22.5 32.5 ;
      RECT 21.5 33.5 22.5 34.5 ;
      RECT 17.5 5.5 18.5 6.5 ;
      RECT 17.5 17.5 18.5 18.5 ;
      RECT 17.5 31.5 18.5 32.5 ;
      RECT 17.5 33.5 18.5 34.5 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 17.5 14.5 18.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 13.5 2.5 14.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END NOR4X1

MACRO OA21X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21X1 0 0 ;
  SIZE 32 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 32 43 ;
        RECT 25 31 27 43 ;
        RECT 21 31 23 43 ;
        RECT 1 31 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 21 13 23 19 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 29 9 31 35 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9 13 11 19 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 17 3 23 ;
    END
  END C
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 32 3 ;
        RECT 25 -3 27 11 ;
        RECT 1 -3 3 11 ;
    END
  END VSS!
  PIN YN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9 21 27 23 ;
        RECT 13 9 19 11 ;
        RECT 13 9 15 23 ;
        RECT 5 31 11 35 ;
        RECT 9 21 11 35 ;
    END
  END YN
  OBS
    LAYER Metal1 ;
      RECT 21 5 23 11 ;
      RECT 5 9 11 11 ;
      RECT 9 5 11 11 ;
      RECT 9 5 23 7 ;
      RECT 13 31 19 35 ;
    LAYER Via1 ;
      RECT 29.5 9.5 30.5 10.5 ;
      RECT 29.5 31.5 30.5 32.5 ;
      RECT 29.5 33.5 30.5 34.5 ;
      RECT 25.5 9.5 26.5 10.5 ;
      RECT 25.5 21.5 26.5 22.5 ;
      RECT 25.5 31.5 26.5 32.5 ;
      RECT 25.5 33.5 26.5 34.5 ;
      RECT 21.5 9.5 22.5 10.5 ;
      RECT 21.5 17.5 22.5 18.5 ;
      RECT 21.5 31.5 22.5 32.5 ;
      RECT 21.5 33.5 22.5 34.5 ;
      RECT 17.5 9.5 18.5 10.5 ;
      RECT 17.5 31.5 18.5 32.5 ;
      RECT 17.5 33.5 18.5 34.5 ;
      RECT 13.5 9.5 14.5 10.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 9.5 10.5 10.5 ;
      RECT 9.5 13.5 10.5 14.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 9.5 6.5 10.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 9.5 2.5 10.5 ;
      RECT 1.5 17.5 2.5 18.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END OA21X1

MACRO OAI21X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21X1 0 0 ;
  SIZE 24 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 24 43 ;
        RECT 21 31 23 43 ;
        RECT 1 31 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 13 3 19 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 13 31 19 35 ;
        RECT 13 21 15 35 ;
        RECT 9 21 15 23 ;
        RECT 9 9 11 23 ;
        RECT 5 9 11 11 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 13 13 15 19 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 21 17 23 23 ;
    END
  END C
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 24 3 ;
        RECT 21 -3 23 11 ;
    END
  END VSS!
  OBS
    LAYER Metal1 ;
      RECT 13 9 19 11 ;
      RECT 1 5 3 11 ;
      RECT 15 5 17 11 ;
      RECT 1 5 17 7 ;
      RECT 5 31 11 35 ;
    LAYER Via1 ;
      RECT 21.5 9.5 22.5 10.5 ;
      RECT 21.5 17.5 22.5 18.5 ;
      RECT 21.5 31.5 22.5 32.5 ;
      RECT 21.5 33.5 22.5 34.5 ;
      RECT 17.5 9.5 18.5 10.5 ;
      RECT 17.5 31.5 18.5 32.5 ;
      RECT 17.5 33.5 18.5 34.5 ;
      RECT 13.5 9.5 14.5 10.5 ;
      RECT 13.5 13.5 14.5 14.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 9.5 10.5 10.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 9.5 6.5 10.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 9.5 2.5 10.5 ;
      RECT 1.5 17.5 2.5 18.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END OAI21X1

MACRO OR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X1 0 0 ;
  SIZE 24 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 24 43 ;
        RECT 17 31 19 43 ;
        RECT 1 31 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 9 3 15 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9 17 11 23 ;
    END
  END B
  PIN YN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 13 21 19 23 ;
        RECT 13 5 15 35 ;
        RECT 5 9 15 11 ;
        RECT 5 5 7 11 ;
    END
  END YN
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 24 3 ;
        RECT 17 -3 19 7 ;
        RECT 9 -3 11 7 ;
        RECT 1 -3 3 7 ;
    END
  END VSS!
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 21 5 23 35 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 5 31 11 35 ;
    LAYER Via1 ;
      RECT 21.5 5.5 22.5 6.5 ;
      RECT 21.5 31.5 22.5 32.5 ;
      RECT 21.5 33.5 22.5 34.5 ;
      RECT 17.5 5.5 18.5 6.5 ;
      RECT 17.5 21.5 18.5 22.5 ;
      RECT 17.5 31.5 18.5 32.5 ;
      RECT 17.5 33.5 18.5 34.5 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 21.5 10.5 22.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 13.5 2.5 14.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END OR2X1

MACRO OR3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3X1 0 0 ;
  SIZE 32 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 32 43 ;
        RECT 25 31 27 43 ;
        RECT 1 31 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 9 3 15 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9 17 11 23 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 17 21 19 27 ;
    END
  END C
  PIN YN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 21 21 27 23 ;
        RECT 21 5 23 35 ;
        RECT 5 9 23 11 ;
        RECT 13 5 15 11 ;
        RECT 5 5 7 11 ;
    END
  END YN
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 32 3 ;
        RECT 25 -3 27 7 ;
        RECT 17 -3 19 7 ;
        RECT 9 -3 11 7 ;
        RECT 1 -3 3 7 ;
    END
  END VSS!
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 29 5 31 35 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 13 31 19 35 ;
      RECT 5 31 11 35 ;
    LAYER Via1 ;
      RECT 29.5 5.5 30.5 6.5 ;
      RECT 29.5 31.5 30.5 32.5 ;
      RECT 29.5 33.5 30.5 34.5 ;
      RECT 25.5 5.5 26.5 6.5 ;
      RECT 25.5 21.5 26.5 22.5 ;
      RECT 25.5 31.5 26.5 32.5 ;
      RECT 25.5 33.5 26.5 34.5 ;
      RECT 21.5 5.5 22.5 6.5 ;
      RECT 21.5 31.5 22.5 32.5 ;
      RECT 21.5 33.5 22.5 34.5 ;
      RECT 17.5 5.5 18.5 6.5 ;
      RECT 17.5 21.5 18.5 22.5 ;
      RECT 17.5 31.5 18.5 32.5 ;
      RECT 17.5 33.5 18.5 34.5 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 21.5 10.5 22.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 13.5 2.5 14.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END OR3X1

MACRO OR4X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4X1 0 0 ;
  SIZE 40 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 40 43 ;
        RECT 33 31 35 43 ;
        RECT 1 31 3 43 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 9 3 15 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9 17 15 19 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 17 17 19 23 ;
    END
  END C
  PIN YN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 29 21 35 23 ;
        RECT 29 5 31 35 ;
        RECT 5 9 31 11 ;
        RECT 21 5 23 11 ;
        RECT 13 5 15 11 ;
        RECT 5 5 7 11 ;
    END
  END YN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 25 21 27 27 ;
    END
  END D
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 40 3 ;
        RECT 33 -3 35 7 ;
        RECT 25 -3 27 7 ;
        RECT 17 -3 19 7 ;
        RECT 9 -3 11 7 ;
        RECT 1 -3 3 7 ;
    END
  END VSS!
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 37 5 39 35 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 21 31 27 35 ;
      RECT 13 31 19 35 ;
      RECT 5 31 11 35 ;
    LAYER Via1 ;
      RECT 37.5 5.5 38.5 6.5 ;
      RECT 37.5 31.5 38.5 32.5 ;
      RECT 37.5 33.5 38.5 34.5 ;
      RECT 33.5 5.5 34.5 6.5 ;
      RECT 33.5 21.5 34.5 22.5 ;
      RECT 33.5 31.5 34.5 32.5 ;
      RECT 33.5 33.5 34.5 34.5 ;
      RECT 29.5 5.5 30.5 6.5 ;
      RECT 29.5 31.5 30.5 32.5 ;
      RECT 29.5 33.5 30.5 34.5 ;
      RECT 25.5 5.5 26.5 6.5 ;
      RECT 25.5 21.5 26.5 22.5 ;
      RECT 25.5 31.5 26.5 32.5 ;
      RECT 25.5 33.5 26.5 34.5 ;
      RECT 21.5 5.5 22.5 6.5 ;
      RECT 21.5 31.5 22.5 32.5 ;
      RECT 21.5 33.5 22.5 34.5 ;
      RECT 17.5 5.5 18.5 6.5 ;
      RECT 17.5 17.5 18.5 18.5 ;
      RECT 17.5 31.5 18.5 32.5 ;
      RECT 17.5 33.5 18.5 34.5 ;
      RECT 13.5 5.5 14.5 6.5 ;
      RECT 13.5 17.5 14.5 18.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 13.5 33.5 14.5 34.5 ;
      RECT 9.5 5.5 10.5 6.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 9.5 33.5 10.5 34.5 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 9.5 2.5 10.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END OR4X1

MACRO TIEHI
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TIEHI 0 0 ;
  SIZE 8 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5 25 7 35 ;
    END
  END Y
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 8 43 ;
        RECT 1 31 3 43 ;
    END
  END VDD!
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 8 3 ;
        RECT 5 -3 7 7 ;
    END
  END VSS!
  OBS
    LAYER Metal1 ;
      RECT 1 5 3 11 ;
    LAYER Via1 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 9.5 2.5 10.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END TIEHI

MACRO TIELO
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TIELO 0 0 ;
  SIZE 8 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5 5 7 11 ;
    END
  END Y
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 8 3 ;
        RECT 1 -3 3 7 ;
    END
  END VSS!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 8 43 ;
        RECT 5 31 7 43 ;
    END
  END VDD!
  OBS
    LAYER Metal1 ;
      RECT 1 25 3 35 ;
    LAYER Via1 ;
      RECT 5.5 5.5 6.5 6.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 5.5 33.5 6.5 34.5 ;
      RECT 1.5 5.5 2.5 6.5 ;
      RECT 1.5 25.5 2.5 26.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
      RECT 1.5 33.5 2.5 34.5 ;
  END
END TIELO

MACRO XNOR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2X1 0 0 ;
  SIZE 40 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 40 3 ;
        RECT 29 -3 31 11 ;
        RECT 17 -3 19 11 ;
        RECT 1 -3 3 11 ;
    END
  END VSS!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 21 3 27 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9 13 11 19 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 33 21 39 23 ;
        RECT 37 9 39 23 ;
        RECT 29 29 35 33 ;
        RECT 33 21 35 33 ;
    END
  END Y
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 40 43 ;
        RECT 37 29 39 43 ;
        RECT 17 29 19 43 ;
        RECT 13 29 15 43 ;
        RECT 1 29 3 43 ;
    END
  END VDD!
  OBS
    LAYER Metal1 ;
      RECT 25 13 35 15 ;
      RECT 33 9 35 15 ;
      RECT 25 9 27 15 ;
      RECT 21 9 27 11 ;
      RECT 5 29 11 33 ;
      RECT 9 21 11 33 ;
      RECT 9 21 15 23 ;
      RECT 13 9 15 23 ;
      RECT 13 17 35 19 ;
      RECT 21 29 27 33 ;
      RECT 5 9 11 11 ;
    LAYER Via1 ;
      RECT 37.5 9.5 38.5 10.5 ;
      RECT 37.5 29.5 38.5 30.5 ;
      RECT 37.5 31.5 38.5 32.5 ;
      RECT 33.5 9.5 34.5 10.5 ;
      RECT 33.5 17.5 34.5 18.5 ;
      RECT 33.5 29.5 34.5 30.5 ;
      RECT 33.5 31.5 34.5 32.5 ;
      RECT 29.5 9.5 30.5 10.5 ;
      RECT 29.5 29.5 30.5 30.5 ;
      RECT 29.5 31.5 30.5 32.5 ;
      RECT 25.5 9.5 26.5 10.5 ;
      RECT 25.5 29.5 26.5 30.5 ;
      RECT 25.5 31.5 26.5 32.5 ;
      RECT 21.5 9.5 22.5 10.5 ;
      RECT 21.5 29.5 22.5 30.5 ;
      RECT 21.5 31.5 22.5 32.5 ;
      RECT 17.5 9.5 18.5 10.5 ;
      RECT 17.5 29.5 18.5 30.5 ;
      RECT 17.5 31.5 18.5 32.5 ;
      RECT 13.5 9.5 14.5 10.5 ;
      RECT 13.5 29.5 14.5 30.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 9.5 9.5 10.5 10.5 ;
      RECT 9.5 13.5 10.5 14.5 ;
      RECT 9.5 29.5 10.5 30.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 5.5 9.5 6.5 10.5 ;
      RECT 5.5 29.5 6.5 30.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 1.5 9.5 2.5 10.5 ;
      RECT 1.5 25.5 2.5 26.5 ;
      RECT 1.5 29.5 2.5 30.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
  END
END XNOR2X1

MACRO XOR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2X1 0 0 ;
  SIZE 40 BY 40 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -3 40 3 ;
        RECT 37 -3 39 11 ;
        RECT 17 -3 19 11 ;
        RECT 13 -3 15 11 ;
        RECT 1 -3 3 11 ;
    END
  END VSS!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 13 3 19 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9 21 11 27 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 37 13 39 33 ;
        RECT 33 13 39 15 ;
        RECT 33 9 35 15 ;
        RECT 29 9 35 11 ;
    END
  END Y
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 37 40 43 ;
        RECT 29 29 31 43 ;
        RECT 17 29 19 43 ;
        RECT 1 29 3 43 ;
    END
  END VDD!
  OBS
    LAYER Metal1 ;
      RECT 13 13 15 33 ;
      RECT 13 17 35 19 ;
      RECT 9 13 15 15 ;
      RECT 9 9 11 15 ;
      RECT 5 9 11 11 ;
      RECT 33 25 35 33 ;
      RECT 21 29 27 33 ;
      RECT 25 25 27 33 ;
      RECT 25 25 35 27 ;
      RECT 21 9 27 11 ;
      RECT 5 29 11 33 ;
    LAYER Via1 ;
      RECT 37.5 9.5 38.5 10.5 ;
      RECT 37.5 29.5 38.5 30.5 ;
      RECT 37.5 31.5 38.5 32.5 ;
      RECT 33.5 9.5 34.5 10.5 ;
      RECT 33.5 17.5 34.5 18.5 ;
      RECT 33.5 29.5 34.5 30.5 ;
      RECT 33.5 31.5 34.5 32.5 ;
      RECT 29.5 9.5 30.5 10.5 ;
      RECT 29.5 29.5 30.5 30.5 ;
      RECT 29.5 31.5 30.5 32.5 ;
      RECT 25.5 9.5 26.5 10.5 ;
      RECT 25.5 29.5 26.5 30.5 ;
      RECT 25.5 31.5 26.5 32.5 ;
      RECT 21.5 9.5 22.5 10.5 ;
      RECT 21.5 29.5 22.5 30.5 ;
      RECT 21.5 31.5 22.5 32.5 ;
      RECT 17.5 9.5 18.5 10.5 ;
      RECT 17.5 29.5 18.5 30.5 ;
      RECT 17.5 31.5 18.5 32.5 ;
      RECT 13.5 9.5 14.5 10.5 ;
      RECT 13.5 29.5 14.5 30.5 ;
      RECT 13.5 31.5 14.5 32.5 ;
      RECT 9.5 9.5 10.5 10.5 ;
      RECT 9.5 25.5 10.5 26.5 ;
      RECT 9.5 29.5 10.5 30.5 ;
      RECT 9.5 31.5 10.5 32.5 ;
      RECT 5.5 9.5 6.5 10.5 ;
      RECT 5.5 29.5 6.5 30.5 ;
      RECT 5.5 31.5 6.5 32.5 ;
      RECT 1.5 9.5 2.5 10.5 ;
      RECT 1.5 13.5 2.5 14.5 ;
      RECT 1.5 29.5 2.5 30.5 ;
      RECT 1.5 31.5 2.5 32.5 ;
  END
END XOR2X1

END LIBRARY
