//Verilog HDL for "KISTA_SOI_STDLIB2", "DECAP4" "functional"


module DECAP4 ( );

endmodule
