*
*
*
*                       LINUX           Thu Dec  2 07:46:02 2021
*
*
*
*  PROGRAM  advgen
*
*  Name           : advgen - Quantus - (64-bit)
*  Version        : 20.1.2-p025
*  Build Date     : Thu Sep 3 13:54:09 PDT 2020
*
*  HSPICE LIBRARY
*
*
*

*
.global VSS! VDD!
.SUBCKT DFFX1 Q D QN CK 
*
*
*  caps2d version: 10
*
*
*       TRANSISTOR CARDS
*
*
MX28_M0_unmatched	QN#2	net055#7	VSS!#1	VSS!#1	nch	L=1e-06
+ W=2e-06
+ AD=5e-12	AS=0	PD=9e-06	PS=0
+ fw=2e-06 sa=2e-06 sb=2e-06
MX27_M0_unmatched	net055#3	qbint#9	VSS!#11	VSS!#11
+ nch	L=1e-06	W=2e-06
+ AD=5e-12	AS=0	PD=9e-06	PS=0	fw=2e-06 sa=2e-06 sb=2e-06
MX26_M0_unmatched	Q#2	qbint#10	VSS!#12	VSS!#12
+ nch	L=1e-06	W=2e-06
+ AD=5e-12	AS=0	PD=9e-06	PS=0	fw=2e-06 sa=2e-06 sb=2e-06
MX25_M0_unmatched	n30#13	CKb#5	net028	net028	nch	L=1e-06
+ W=2e-06
+ AD=5e-12	AS=0	PD=9e-06	PS=0
+ fw=2e-06 sa=2e-06 sb=2e-06
MX24_M0_unmatched	net028#2	qbint#12	VSS!#13	VSS!#13
+ nch	L=1e-06	W=2e-06
+ AD=5e-12	AS=0	PD=9e-06	PS=0	fw=2e-06 sa=2e-06 sb=2e-06
MX23_M0_unmatched	qbint#3	n30#9	VSS!#14	VSS!#14
+ nch	L=1e-06	W=2e-06
+ AD=5e-12	AS=0	PD=9e-06	PS=0	fw=2e-06 sa=2e-06 sb=2e-06
MX22_M0_unmatched	n30#4	CKbb#9	mout#11	mout#11	nch
+ L=1e-06	W=2e-06
+ AD=5e-12	AS=0	PD=9e-06	PS=0
+ fw=2e-06 sa=2e-06 sb=2e-06
MX21_M0_unmatched	n20#12	CKbb#10	net017	net017	nch	L=1e-06
+ W=2e-06
+ AD=5e-12	AS=0	PD=9e-06	PS=0
+ fw=2e-06 sa=2e-06 sb=2e-06
MX20_M0_unmatched	net017#2	mout#4	VSS!#15	VSS!#15
+ nch	L=1e-06	W=2e-06
+ AD=5e-12	AS=0	PD=9e-06	PS=0	fw=2e-06 sa=2e-06 sb=2e-06
MX19_M0_unmatched	mout#7	n20#8	VSS!#16	VSS!#16	nch
+ L=1e-06	W=2e-06
+ AD=5e-12	AS=0	PD=9e-06	PS=0
+ fw=2e-06 sa=2e-06 sb=2e-06
MX18_M0_unmatched	n20#3	CKb#13	net13	net13	nch	L=1e-06
+ W=2e-06
+ AD=5e-12	AS=0	PD=9e-06	PS=0
+ fw=2e-06 sa=2e-06 sb=2e-06
MX17_M0_unmatched	net13#2	D#3	VSS!#17	VSS!#17
+ nch	L=1e-06	W=2e-06
+ AD=5e-12	AS=0	PD=9e-06	PS=0	fw=2e-06 sa=2e-06 sb=2e-06
MX16_M0_unmatched	CKbb#4	CKb#9	VSS!#18	VSS!#18	nch
+ L=1e-06	W=2e-06
+ AD=5e-12	AS=0	PD=9e-06	PS=0
+ fw=2e-06 sa=2e-06 sb=2e-06
MX15_M0_unmatched	CKb#3	CK#4	VSS!#10	VSS!#10	nch
+ L=1e-06	W=2e-06
+ AD=5e-12	AS=0	PD=9e-06	PS=0
+ fw=2e-06 sa=2e-06 sb=2e-06
MX42_M0_unmatched	QN#3	net055#5	VDD!#1	VDD!#1	pch	L=1e-06
+ W=4e-06
+ AD=1e-11	AS=0	PD=1.3e-05	PS=0
+ fw=4e-06 sa=2e-06 sb=2e-06
MX41_M0_unmatched	net055#4	qbint#5	VDD!#11	VDD!#11
+ pch	L=1e-06	W=4e-06
+ AD=1e-11	AS=0	PD=1.3e-05	PS=0	fw=4e-06 sa=2e-06 sb=2e-06
MX40_M0_unmatched	Q#3	qbint#11	VDD!#12	VDD!#12
+ pch	L=1e-06	W=4e-06
+ AD=1e-11	AS=0	PD=1.3e-05	PS=0	fw=4e-06 sa=2e-06 sb=2e-06
MX39_M0_unmatched	n30#10	CKbb#5	net029	net029	pch	L=1e-06
+ W=4e-06
+ AD=1e-11	AS=0	PD=1.3e-05	PS=0
+ fw=4e-06 sa=2e-06 sb=2e-06
MX38_M0_unmatched	net029#2	qbint#13	VDD!#13	VDD!#13
+ pch	L=1e-06	W=4e-06
+ AD=1e-11	AS=0	PD=1.3e-05	PS=0	fw=4e-06 sa=2e-06 sb=2e-06
MX37_M0_unmatched	qbint#4	n30#7	VDD!#14	VDD!#14
+ pch	L=1e-06	W=4e-06
+ AD=1e-11	AS=0	PD=1.3e-05	PS=0	fw=4e-06 sa=2e-06 sb=2e-06
MX36_M0_unmatched	n30#5	CKb#11	mout#9	mout#9	pch	L=1e-06
+ W=4e-06
+ AD=1e-11	AS=0	PD=1.3e-05	PS=0
+ fw=4e-06 sa=2e-06 sb=2e-06
MX35_M0_unmatched	n20#10	CKb#12	net018	net018	pch	L=1e-06
+ W=4e-06
+ AD=1e-11	AS=0	PD=1.3e-05	PS=0
+ fw=4e-06 sa=2e-06 sb=2e-06
MX34_M0_unmatched	net018#2	mout	VDD!#15	VDD!#15
+ pch	L=1e-06	W=4e-06
+ AD=1e-11	AS=0	PD=1.3e-05	PS=0	fw=4e-06 sa=2e-06 sb=2e-06
MX33_M0_unmatched	mout#8	n20#6	VDD!#16	VDD!#16	pch
+ L=1e-06	W=4e-06
+ AD=1e-11	AS=0	PD=1.3e-05	PS=0
+ fw=4e-06 sa=2e-06 sb=2e-06
MX32_M0_unmatched	n20#5	CKbb#11	net14	net14	pch	L=1e-06
+ W=4e-06
+ AD=1e-11	AS=0	PD=1.3e-05	PS=0
+ fw=4e-06 sa=2e-06 sb=2e-06
MX31_M0_unmatched	net14#2	D#2	VDD!#17	VDD!#17
+ pch	L=1e-06	W=4e-06
+ AD=1e-11	AS=0	PD=1.3e-05	PS=0	fw=4e-06 sa=2e-06 sb=2e-06
MX30_M0_unmatched	CKbb#2	CKb#14	VDD!#18	VDD!#18	pch
+ L=1e-06	W=4e-06
+ AD=1e-11	AS=0	PD=1.3e-05	PS=0
+ fw=4e-06 sa=2e-06 sb=2e-06
MX29_M0_unmatched	CKb#4	CK#2	VDD!#10	VDD!#10	pch
+ L=1e-06	W=4e-06
+ AD=1e-11	AS=0	PD=1.3e-05	PS=0
+ fw=4e-06 sa=2e-06 sb=2e-06
*
*
*       RESISTOR AND CAP/DIODE CARDS
*
Rd4	D#2	D#1	  927.2892	$poly_conn
Rd5	D#1	D#3	 1347.2892	$poly_conn
Rd28	CKb#6	CKb#11	 3766.2549
Rd22	CKb#7	CKb#12	 3766.2549
Rd29	CKb#8	CKb#9	 2928.0679
Rd23	CKb#10	CKb	   42.9640
Rd30	CKb	CKb#3	   20.2150
Rd25	qbint#5	qbint#6	 1014.2584
Rd24	qbint#6	qbint#7	 1117.6837
Rd31	qbint#7	qbint#10	 1419.0477
Rd26	qbint#8	qbint#13	  997.5659
Rd27	qbint#8	qbint	   82.8419
Rd32	qbint	qbint#3	   20.2150
Rd36	CKbb#5	CKbb#6	 3408.0676
Rd38	CKbb#6	CKbb#7	 1188.5167
Rd37	CKbb#7	CKbb#8	 4188.5166
Rd33	CKbb#8	CKbb	 2001.5475
Rd40	CKbb	CKbb#4	   21.8702
Rd39	net055#5	net055#6	 1014.2584
Rd35	net055#6	net055	  445.9252
Rd34	net055	net055#3	   20.0314
Rd12	CK#2	CK#3	 1014.2584
Rd14	CK#3	CK	  450.9377
Rd13	VSS!#1	VSS!#11	  151.6630
Rd15	VSS!#1	VSS!#3	    5.7608
Rd19	VSS!#3	VSS!#13	   15.9906
Rd20	VSS!#13	VSS!#5	    7.9180
Rd16	VSS!#5	VSS!#6	    0.5962
Rd21	VSS!#6	VSS!#16	    7.9180
Rd18	VSS!#6	VSS!#8	    0.6074
Rd17	VSS!#8	VSS!#17	    5.1645
Rd6	VSS!#8	VSS!#18	   10.2888
Rd8	VDD!#1	VDD!#2	    2.9060
Rd7	VDD!#2	VDD!#12	    4.2474
Rd9	VDD!#12	VDD!#4	    8.5777
Rd11	VDD!#4	VDD!#14	    3.7973
Rd10	VDD!#14	VDD!#6	   11.5401
Rd41	VDD!#6	VDD!#16	    4.2474
Rd43	VDD!#6	VDD!#8	    0.6210
Rd42	VDD!#8	VDD!#17	    2.7095
Rd1	VDD!#8	VDD!#18	    5.5891
Rd3	n30#8	n30#9	 1426.0319
Rd2	n30	n30#2	    5.0795
Rc8	D	D#1	    5.0025	$metal1_conn
Rc41	Q	Q#3	    2.7206	$metal1_conn
Rc40	Q	Q#2	    5.2606	$metal1_conn
Rc47	QN	QN#3	    2.8181	$metal1_conn
Rc46	QN	QN#2	    5.1631	$metal1_conn
Rc15	net018	net018#2	    5.0750	$metal1_conn
Rc34	net029	net029#2	    5.0750	$metal1_conn
Rc9	net14	net14#2	    5.0750	$metal1_conn
Rc35	net028	net028#2	   10.1000	$metal1_conn
Rc10	net13	net13#2	   10.1000	$metal1_conn
Rc16	net017	net017#2	   10.1000	$metal1_conn
Rc75	CKb#6	CKb#5	 4728.0679
Rc66	CKb#7	CKb#8	 2988.5168
Rc76	CKb#9	CKb#10	 1426.0319
Rc77	CKb	CKb#4	   10.4399
Rc67	CKb#4	CKb#3	   10.7906
Rc78	qbint#6	qbint#9	 1434.2584
Rc68	qbint#7	qbint#11	  999.0477
Rc79	qbint#7	qbint#8	 2362.7004
Rc69	qbint#8	qbint#12	 1417.5659
Rc80	qbint	qbint#4	   10.4399
Rc70	qbint#4	qbint#3	   10.7906
Rc81	CKbb#6	CKbb#9	 3813.8738
Rc71	CKbb#7	CKbb#10	 3946.2549
Rc82	CKbb#8	CKbb#11	  418.6361
Rc72	CKbb	CKbb#2	    9.9682
Rc74	CKbb#2	CKbb#4	   10.6580
Rc83	net055#6	net055#7	 1434.2584
Rc73	net055	net055#4	   10.3451
Rc57	net055#4	net055#3	   10.8255
Rc48	CK#3	CK#4	 1434.2584
Rc58	VSS!	VSS!#10	    5.1886
Rc59	VSS!#11	VSS!#3	    5.5497
Rc49	VSS!#3	VSS!#12	    5.1645
Rc60	VSS!#3	VSS!#5	    0.6074
Rc50	VSS!#5	VSS!#14	    5.1645
Rc61	VSS!#6	VSS!#15	    5.1645
Rc51	VSS!	VSS!#8	    0.4096
Rc62	VSS!#16	VSS!#8	   15.9906
Rc52	VSS!	VSS!#18	   10.7825
Rc63	VDD!	VDD!#10	    2.7386
Rc53	VDD!#2	VDD!#11	    2.7095
Rc64	VDD!#2	VDD!#4	    0.6210
Rc54	VDD!#4	VDD!#13	    2.7095
Rc56	VDD!#4	VDD!#6	    0.8355
Rc65	VDD!#6	VDD!#15	    2.7095
Rc55	VDD!	VDD!#8	    0.4086
Rc2	VDD!#16	VDD!#8	    8.5777
Rc4	VDD!	VDD!#18	    5.6436
Rc3	n30#7	n30#8	 1006.0318
Rc31	n30#8	n30	   80.4640
Rc33	n30#2	n30#5	    2.7181
Rc32	n30#2	n30#4	    5.1631
Rc26	n30#2	n30#10	    3.9915
Rc30	n30#2	n30#13	    7.3129
Rc29	n30#10	n30#13	   27.1489
Rc28	n20#6	n20#7	 1014.2584
Rc37	n20#7	n20#8	 1434.2584
Rc36	n20#7	n20#2	  750.9252
Rc38	n20#2	n20	    0.1745
Rc5	n20#2	n20#5	    2.7200
Rc7	n20#2	n20#3	    5.1631
Rc6	n20	n20#10	    3.7217
Rc11	n20	n20#12	    6.8186
Rc14	n20#10	n20#12	   32.8723
Rc12	mout	mout#2	 1006.0318
Rc22	mout#2	mout#4	 1426.0319
Rc21	mout#2	mout#3	   47.9640
Rc23	mout#3	mout#9	    3.6110
Rc17	mout#3	mout#11	    6.9897
Rc24	mout#9	mout#11	   32.3608
Rc25	mout#3	mout#8	    2.7181
Rc20	mout#3	mout#7	    5.2631
Rb3	CKb#6	CKb#7	 1188.5167
Rb1	CKb#8	CKb#13	  538.6361
Rb2	CKb#10	CKb#14	 1006.0318
*
*       CAPACITOR CARDS
*
*
C1	VSS!	Q	2.98659e-15
C2	Q#3	VSS!	9.51892e-16
C3	Q#2	VSS!	1.14529e-15
C4	VSS!	D	3.51676e-16
C5	D#2	VSS!	1.81618e-15
C6	D#3	VSS!	2.17032e-15
C7	D#1	VSS!	3.75027e-15
C8	VSS!	QN	2.99091e-15
C9	QN#3	VSS!	1.77117e-15
C10	QN#2	VSS!	8.80953e-16
C11	VSS!	CK	1.94402e-15
C12	CK#2	VSS!	1.94399e-15
C13	CK#4	VSS!	2.37844e-15
C14	CK#3	VSS!	3.45207e-15
C15	VDD!	VSS!	6.93391e-17
C16	VDD!#1	VSS!	5.06526e-16
C17	VDD!#11	VSS!	4.76565e-16
C18	VDD!#12	VSS!	4.96774e-16
C19	VDD!#13	VSS!	1.1943e-15
C20	VDD!#14	VSS!	1.05168e-15
C21	VDD!#15	VSS!	8.68992e-16
C22	VDD!#16	VSS!	7.78974e-16
C23	VDD!#17	VSS!	8.23361e-16
C24	VDD!#18	VSS!	5.86659e-16
C25	VDD!#10	VSS!	6.73761e-16
C26	VDD!#6	VSS!	2.87597e-15
C27	CKb#11	VSS!	1.86429e-15
C28	CKb#12	VSS!	1.81604e-15
C29	CKb#14	VSS!	9.55665e-16
C30	CKb#5	VSS!	1.18287e-15
C31	CKb#13	VSS!	2.48461e-16
C32	CKb#9	VSS!	1.0494e-15
C33	CKb#4	VSS!	2.09801e-15
C34	CKb#6	VSS!	1.65962e-15
C35	CKb#7	VSS!	2.06769e-15
C36	CKb#8	VSS!	1.28355e-15
C37	CKbb#5	VSS!	1.0804e-15
C38	CKbb#11	VSS!	9.07339e-16
C39	CKbb#9	VSS!	2.4533e-15
C40	CKbb#10	VSS!	1.67105e-15
C41	CKbb#2	VSS!	2.42466e-15
C42	CKbb#6	VSS!	3.52021e-15
C43	CKbb#7	VSS!	2.3095e-15
C44	CKbb#8	VSS!	1.17949e-15
C45	n20	VSS!	7.16217e-15
C46	n20#6	VSS!	9.59367e-16
C47	n20#8	VSS!	3.52428e-16
C48	n20#7	VSS!	2.41586e-16
C49	mout	VSS!	8.54558e-16
C50	mout#4	VSS!	2.32808e-16
C51	mout#3	VSS!	7.15315e-15
C52	n30#7	VSS!	9.65203e-16
C53	n30#9	VSS!	3.56919e-16
C54	n30#2	VSS!	8.23852e-15
C55	qbint#5	VSS!	9.6256e-16
C56	qbint#11	VSS!	9.62419e-16
C57	qbint#13	VSS!	8.45216e-16
C58	qbint#9	VSS!	3.76151e-16
C59	qbint#10	VSS!	3.76011e-16
C60	qbint#12	VSS!	2.33255e-16
C61	qbint#4	VSS!	2.93652e-15
C62	qbint#6	VSS!	6.09929e-16
C63	qbint#7	VSS!	1.64578e-15
C64	net055#5	VSS!	9.21882e-16
C65	net055#7	VSS!	3.57581e-16
C66	net055#4	VSS!	1.27654e-15
C67	net055#6	VSS!	2.82077e-16
C68	VSS!	VSS!	6.4805e-14
C69	net13	VSS!	3.8404e-16
C70	net13#2	VSS!	4.20384e-16
C71	net017	VSS!	5.8867e-16
C72	net017#2	VSS!	5.75009e-16
C73	net028	VSS!	4.02281e-16
C74	net028#2	VSS!	4.15914e-16
C75	net14	VSS!	4.80482e-16
C76	net14#2	VSS!	5.16663e-16
C77	net018	VSS!	4.68993e-16
C78	net018#2	VSS!	4.62138e-16
C79	net029	VSS!	5.50503e-16
C80	net029#2	VSS!	5.65584e-16
C81	X42_5	VSS!	1.14629e-15
C82	X41_5	VSS!	8.79514e-16
C83	X40_5	VSS!	8.42637e-16
C84	X39_5	VSS!	8.9421e-16
C85	X38_5	VSS!	9.43004e-16
C86	X37_5	VSS!	1.49843e-15
C87	X36_5	VSS!	1.89839e-15
C88	X35_5	VSS!	1.38155e-15
C89	X34_5	VSS!	9.57117e-16
C90	X33_5	VSS!	9.54453e-16
C91	X32_5	VSS!	9.39862e-16
C92	X31_5	VSS!	8.70159e-16
C93	X30_5	VSS!	1.0676e-15
C94	X29_5	VSS!	1.1697e-15
C95	VDD!#2	VSS!	4.03266e-14
C96	VSS!	CKb	4.36954e-15
C97	CKb#11	VSS!	3.96668e-15
C98	CKb#12	VSS!	4.52014e-15
C99	CKb#14	VSS!	8.94338e-16
C100	CKb#5	VSS!	5.88243e-15
C101	CKb#13	VSS!	1.42424e-15
C102	CKb#9	VSS!	4.58728e-15
C103	CKb#4	VSS!	2.19835e-15
C104	CKb#3	VSS!	9.76506e-16
C105	CKb#6	VSS!	9.85802e-15
C106	CKb#7	VSS!	7.9493e-15
C107	CKb#8	VSS!	6.34425e-15
C108	VSS!	CKbb	3.57961e-15
C109	CKbb#5	VSS!	4.16052e-15
C110	CKbb#11	VSS!	7.31822e-16
C111	CKbb#9	VSS!	4.61267e-15
C112	CKbb#10	VSS!	4.95155e-15
C113	CKbb#2	VSS!	1.47931e-15
C114	CKbb#4	VSS!	1.65854e-15
C115	CKbb#6	VSS!	7.62996e-15
C116	CKbb#7	VSS!	8.28618e-15
C117	CKbb#8	VSS!	6.74423e-15
C118	n20#6	VSS!	1.00187e-15
C119	n20#8	VSS!	1.98471e-15
C120	n20#2	VSS!	1.04885e-14
C121	n20#7	VSS!	3.44683e-15
C122	VSS!	mout	9.16272e-16
C123	mout#4	VSS!	1.93316e-15
C124	mout#3	VSS!	1.14346e-14
C125	n30#7	VSS!	8.86643e-16
C126	n30#9	VSS!	1.88667e-15
C127	n30#2	VSS!	1.24046e-14
C128	VSS!	qbint	6.82682e-15
C129	qbint#5	VSS!	9.91231e-16
C130	qbint#11	VSS!	9.91562e-16
C131	qbint#13	VSS!	9.26825e-16
C132	qbint#9	VSS!	2.01378e-15
C133	qbint#10	VSS!	2.01378e-15
C134	qbint#12	VSS!	1.92327e-15
C135	qbint#4	VSS!	2.38123e-15
C136	qbint#3	VSS!	8.70725e-16
C137	qbint#6	VSS!	3.80757e-15
C138	qbint#7	VSS!	6.03785e-15
C139	VSS!	net055	1.63853e-15
C140	net055#5	VSS!	9.7896e-16
C141	net055#7	VSS!	1.97197e-15
C142	net055#4	VSS!	2.15147e-15
C143	net055#3	VSS!	8.00821e-16
C144	net055#6	VSS!	3.10866e-15
*
*
.ENDS DFFX1
*
