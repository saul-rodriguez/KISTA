//Verilog HDL for "KISTA_SOI_STDLIB2", "DECAP3" "functional"


module DECAP3 ( );

endmodule
