*
*
*
*                       LINUX           Tue Dec 21 06:03:40 2021
*
*
*
*  PROGRAM  advgen
*
*  Name           : advgen - Quantus - (64-bit)
*  Version        : 20.1.2-p025
*  Build Date     : Thu Sep 3 13:54:09 PDT 2020
*
*  HSPICE LIBRARY
*
*
*

*
.GLOBAL VSS! VDD!
.SUBCKT AOI21X1 A0 Y B0 A1
*
*
*  caps2d version: 10
*
*
*       TRANSISTOR CARDS
*
*
MX8_M0_unmatched	Y#3	B0#4	VSS!#2	VSS!#2	nch	L=1e-06
+ W=2e-06
+ AD=5e-12	AS=0	PD=9e-06	PS=0
+ fw=2e-06 sa=2e-06 sb=2e-06
MX4_M0_unmatched	Y#4	A0#4	net17	net17	nch	L=1e-06
+ W=4e-06
+ AD=1e-11	AS=0	PD=1.3e-05	PS=0
+ fw=4e-06 sa=2e-06 sb=2e-06
MX3_M0_unmatched	net17#2	A1#6	VSS!#1	VSS!#1	nch	L=1e-06
+ W=4e-06
+ AD=1e-11	AS=0	PD=1.3e-05	PS=0
+ fw=4e-06 sa=2e-06 sb=2e-06
MX7_M0_unmatched	Y#1	A0#2	net19	net19	pch	L=1e-06
+ W=8e-06
+ AD=2e-11	AS=0	PD=2.1e-05	PS=0
+ fw=8e-06 sa=2e-06 sb=2e-06
MX6_M0_unmatched	Y#5	A1#4	net19#4	net19#4	pch
+ L=1e-06	W=8e-06
+ AD=2e-11	AS=0	PD=2.1e-05	PS=0
+ fw=8e-06 sa=2e-06 sb=2e-06
MX5_M0_unmatched	net19#3	B0#2	VDD!#1	VDD!#1	pch	L=1e-06
+ W=8e-06
+ AD=2e-11	AS=0	PD=2.1e-05	PS=0
+ fw=8e-06 sa=2e-06 sb=2e-06
*
*
*       RESISTOR AND CAP/DIODE CARDS
*
Rd4	A1#4	A1#5	  957.2891
Rd5	A1#5	A1	    5.0512
Rd6	Y	Y#4	    2.8150
Rd7	Y#5	Y#3	   32.1847
Rd9	A0#2	A0#3	 1636.0317
Rd8	A0#3	A0	   85.4690
Rd1	B0#3	B0#4	 1936.0317
Rd3	net19	net19#4	    3.7950
Rd2	net19#4	net19#3	    4.6089
Rc15	VSS!#1	VSS!	    2.6779	$metal1_conn
Rc16	VSS!	VSS!#2	    5.2044	$metal1_conn
Rc9	net17	net17#2	    5.0750	$metal1_conn
Rc17	VDD!	VDD!#1	    1.5694	$metal1_conn
Rc2	A1#5	A1#6	  957.2891
Rc3	Y#1	Y	    1.4350
Rc4	Y	Y#5	    1.7829
Rc10	Y	Y#3	    6.8878
Rc13	A0#3	A0#4	  436.0318
Rc11	B0#2	B0#3	  436.0318
Rc14	B0#3	B0	   85.4690
Rc12	net19	net19#3	    4.8158
Rs1		4	VSS!	50
*
*       CAPACITOR CARDS
*
*
C1	Y	A0	1.42714e-16
C2	A0#2	Y	8.572e-16
C3	Y#4	A0	1.82029e-16
C4	Y#4	A0#4	1.56192e-16
C5	A0#3	Y	1.66163e-17
C6	VSS!	A0	1.16358e-17
C7	A0#2	VSS!	6.37688e-18
C8	A0#4	VSS!	6.54153e-17
C9	A0#3	VSS!	1.19556e-19
C10	A0#2	VDD!	1.09299e-17
C11	A1	A0	4.03514e-18
C12	A1#5	A0	4.13602e-20
C13	A0#3	A1	2.50993e-19
C14	A0#3	A1#5	2.57267e-21
C15	4	A0	3.80431e-15
C16	A0#2	4	1.49001e-15
C17	A0#4	4	7.82769e-16
C18	A0#3	4	2.24262e-16
C19	net17	A0	5.06958e-17
C20	A0#4	net17	1.3805e-16
C21	A0#3	net17	7.3974e-19
C22	A0#2	net19	2.47754e-16
C23	A0#2	X7_5	5.0433e-16
C24	B0	Y	2.93557e-16
C25	Y#3	B0	3.45358e-17
C26	Y#3	B0#4	2.74546e-16
C27	Y#4	VSS!	8.76192e-17
C28	Y#3	VSS!#1	1.68727e-16
C29	Y#1	VDD!	1.39618e-17
C30	A1	Y	4.18236e-16
C31	Y#5	A1#4	5.77632e-16
C32	Y#3	A1	5.78523e-18
C33	Y#3	A1#6	1.13428e-17
C34	A1#5	Y	3.48892e-18
C35	4	Y	5.98803e-15
C36	Y#1	4	5.67488e-17
C37	Y#4	4	1.48327e-15
C38	Y#5	4	5.61811e-17
C39	Y#3	4	1.5977e-15
C40	Y#4	net17	7.91422e-17
C41	net17#2	Y	3.62116e-18
C42	net19	Y	5.25258e-17
C43	Y#1	net19	1.40494e-16
C44	net19#4	Y	5.80138e-17
C45	net19#3	Y	5.18397e-17
C46	net19#3	Y#5	2.73208e-16
C47	Y#1	X7_5	6.46972e-16
C48	Y#5	X6_5	2.26143e-16
C49	VSS!	B0	4.5743e-18
C50	B0#2	VSS!	1.08435e-17
C51	VSS!#2	B0	2.29042e-18
C52	VSS!#2	B0#4	1.90428e-16
C53	VDD!#1	B0	5.34874e-17
C54	VDD!#1	B0#2	2.89384e-16
C55	4	B0	4.37052e-15
C56	B0#2	4	2.93574e-16
C57	B0#4	4	2.46027e-15
C58	B0#3	4	2.43142e-19
C59	net19#3	B0#2	2.76012e-16
C60	B0#2	X5_5	5.32553e-16
C61	VDD!	VSS!	7.32018e-18
C62	A1	VSS!	9.0072e-18
C63	A1#4	VSS!	1.39104e-17
C64	VSS!#1	A1	7.48118e-18
C65	VSS!#1	A1#6	2.42912e-16
C66	4	VSS!	4.91368e-15
C67	VSS!#1	4	5.28518e-16
C68	VSS!#2	4	1.84609e-15
C69	net17	VSS!	7.40211e-17
C70	net17#2	VSS!	6.36502e-17
C71	VSS!#1	net17#2	7.21635e-17
C72	net19#4	VSS!	1.17783e-17
C73	4	VDD!	6.76683e-15
C74	VDD!#1	4	7.20267e-16
C75	net19#4	VDD!	2.34304e-16
C76	net19#3	VDD!#1	2.0956e-16
C77	X5_5	VDD!	2.866e-17
C78	VDD!#1	X5_5	6.03838e-16
C79	4	A1	3.73767e-15
C80	A1#4	4	8.57837e-16
C81	A1#6	4	1.42508e-15
C82	A1#5	4	3.28518e-17
C83	net17#2	A1#6	1.38973e-16
C84	net19#4	A1#4	3.53084e-16
C85	A1#4	X6_5	5.10168e-16
C86	net17	4	2.28442e-16
C87	net17#2	4	2.28694e-16
C88	net19#4	4	1.57237e-15
C89	net19#3	4	1.41651e-15
C90	X7_5	net19	1.0929e-16
C91	net19#4	X7_5	7.9165e-17
C92	net19#4	X6_5	3.29742e-16
C93	net19#3	X5_5	1.49036e-16
*
*
.ENDS AOI21X1
*
